VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_0rw1r1w_23_32_freepdk45
   CLASS BLOCK ;
   SIZE 97.4 BY 92.89 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  21.8175 0.0 21.9575 0.14 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  24.6775 0.0 24.8175 0.14 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  27.5375 0.0 27.6775 0.14 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  30.3975 0.0 30.5375 0.14 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  33.2575 0.0 33.3975 0.14 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  36.1175 0.0 36.2575 0.14 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  38.9775 0.0 39.1175 0.14 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  41.8375 0.0 41.9775 0.14 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  44.6975 0.0 44.8375 0.14 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  47.5575 0.0 47.6975 0.14 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  50.4175 0.0 50.5575 0.14 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  53.2775 0.0 53.4175 0.14 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  56.1375 0.0 56.2775 0.14 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  58.9975 0.0 59.1375 0.14 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  61.8575 0.0 61.9975 0.14 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  64.7175 0.0 64.8575 0.14 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  67.5775 0.0 67.7175 0.14 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  70.4375 0.0 70.5775 0.14 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  73.2975 0.0 73.4375 0.14 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  76.1575 0.0 76.2975 0.14 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  79.0175 0.0 79.1575 0.14 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  81.8775 0.0 82.0175 0.14 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  84.7375 0.0 84.8775 0.14 ;
      END
   END din0[22]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 45.815 0.14 45.955 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 48.545 0.14 48.685 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 50.755 0.14 50.895 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 53.485 0.14 53.625 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 55.695 0.14 55.835 ;
      END
   END addr0[4]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.26 22.675 97.4 22.815 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.26 19.945 97.4 20.085 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.26 17.735 97.4 17.875 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  80.835 0.0 80.975 0.14 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  81.12 0.0 81.26 0.14 ;
      END
   END addr1[4]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 4.215 0.14 4.355 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.26 88.535 97.4 88.675 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  9.56 0.0 9.7 0.14 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  87.7 92.75 87.84 92.89 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  35.0475 92.75 35.1875 92.89 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  36.2225 92.75 36.3625 92.89 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  37.3975 92.75 37.5375 92.89 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  38.5725 92.75 38.7125 92.89 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  39.7475 92.75 39.8875 92.89 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  40.9225 92.75 41.0625 92.89 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  42.0975 92.75 42.2375 92.89 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  43.2725 92.75 43.4125 92.89 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  44.4475 92.75 44.5875 92.89 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  45.6225 92.75 45.7625 92.89 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  46.7975 92.75 46.9375 92.89 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  47.9725 92.75 48.1125 92.89 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  49.1475 92.75 49.2875 92.89 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  50.3225 92.75 50.4625 92.89 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  51.4975 92.75 51.6375 92.89 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  52.6725 92.75 52.8125 92.89 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  53.8475 92.75 53.9875 92.89 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  55.0225 92.75 55.1625 92.89 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  56.1975 92.75 56.3375 92.89 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  57.3725 92.75 57.5125 92.89 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  58.5475 92.75 58.6875 92.89 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  59.7225 92.75 59.8625 92.89 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  60.8975 92.75 61.0375 92.89 ;
      END
   END dout1[22]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 97.26 92.75 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 97.26 92.75 ;
   LAYER  metal3 ;
      RECT  0.28 45.675 97.26 46.095 ;
      RECT  0.14 46.095 0.28 48.405 ;
      RECT  0.14 48.825 0.28 50.615 ;
      RECT  0.14 51.035 0.28 53.345 ;
      RECT  0.14 53.765 0.28 55.555 ;
      RECT  0.14 55.975 0.28 92.75 ;
      RECT  0.28 0.14 97.12 22.535 ;
      RECT  0.28 22.535 97.12 22.955 ;
      RECT  0.28 22.955 97.12 45.675 ;
      RECT  97.12 22.955 97.26 45.675 ;
      RECT  97.12 20.225 97.26 22.535 ;
      RECT  97.12 0.14 97.26 17.595 ;
      RECT  97.12 18.015 97.26 19.805 ;
      RECT  0.14 0.14 0.28 4.075 ;
      RECT  0.14 4.495 0.28 45.675 ;
      RECT  0.28 46.095 97.12 88.395 ;
      RECT  0.28 88.395 97.12 88.815 ;
      RECT  0.28 88.815 97.12 92.75 ;
      RECT  97.12 46.095 97.26 88.395 ;
      RECT  97.12 88.815 97.26 92.75 ;
   LAYER  metal4 ;
      RECT  0.14 0.42 21.5375 92.75 ;
      RECT  21.5375 0.42 22.2375 92.75 ;
      RECT  22.2375 0.14 24.3975 0.42 ;
      RECT  25.0975 0.14 27.2575 0.42 ;
      RECT  27.9575 0.14 30.1175 0.42 ;
      RECT  30.8175 0.14 32.9775 0.42 ;
      RECT  33.6775 0.14 35.8375 0.42 ;
      RECT  36.5375 0.14 38.6975 0.42 ;
      RECT  39.3975 0.14 41.5575 0.42 ;
      RECT  42.2575 0.14 44.4175 0.42 ;
      RECT  45.1175 0.14 47.2775 0.42 ;
      RECT  47.9775 0.14 50.1375 0.42 ;
      RECT  50.8375 0.14 52.9975 0.42 ;
      RECT  53.6975 0.14 55.8575 0.42 ;
      RECT  56.5575 0.14 58.7175 0.42 ;
      RECT  59.4175 0.14 61.5775 0.42 ;
      RECT  62.2775 0.14 64.4375 0.42 ;
      RECT  65.1375 0.14 67.2975 0.42 ;
      RECT  67.9975 0.14 70.1575 0.42 ;
      RECT  70.8575 0.14 73.0175 0.42 ;
      RECT  73.7175 0.14 75.8775 0.42 ;
      RECT  76.5775 0.14 78.7375 0.42 ;
      RECT  82.2975 0.14 84.4575 0.42 ;
      RECT  85.1575 0.14 97.26 0.42 ;
      RECT  79.4375 0.14 80.555 0.42 ;
      RECT  81.54 0.14 81.5975 0.42 ;
      RECT  0.14 0.14 9.28 0.42 ;
      RECT  9.98 0.14 21.5375 0.42 ;
      RECT  22.2375 0.42 87.42 92.47 ;
      RECT  87.42 0.42 88.12 92.47 ;
      RECT  88.12 0.42 97.26 92.47 ;
      RECT  88.12 92.47 97.26 92.75 ;
      RECT  22.2375 92.47 34.7675 92.75 ;
      RECT  35.4675 92.47 35.9425 92.75 ;
      RECT  36.6425 92.47 37.1175 92.75 ;
      RECT  37.8175 92.47 38.2925 92.75 ;
      RECT  38.9925 92.47 39.4675 92.75 ;
      RECT  40.1675 92.47 40.6425 92.75 ;
      RECT  41.3425 92.47 41.8175 92.75 ;
      RECT  42.5175 92.47 42.9925 92.75 ;
      RECT  43.6925 92.47 44.1675 92.75 ;
      RECT  44.8675 92.47 45.3425 92.75 ;
      RECT  46.0425 92.47 46.5175 92.75 ;
      RECT  47.2175 92.47 47.6925 92.75 ;
      RECT  48.3925 92.47 48.8675 92.75 ;
      RECT  49.5675 92.47 50.0425 92.75 ;
      RECT  50.7425 92.47 51.2175 92.75 ;
      RECT  51.9175 92.47 52.3925 92.75 ;
      RECT  53.0925 92.47 53.5675 92.75 ;
      RECT  54.2675 92.47 54.7425 92.75 ;
      RECT  55.4425 92.47 55.9175 92.75 ;
      RECT  56.6175 92.47 57.0925 92.75 ;
      RECT  57.7925 92.47 58.2675 92.75 ;
      RECT  58.9675 92.47 59.4425 92.75 ;
      RECT  60.1425 92.47 60.6175 92.75 ;
      RECT  61.3175 92.47 87.42 92.75 ;
   END
END    sram_0rw1r1w_23_32_freepdk45
END    LIBRARY
