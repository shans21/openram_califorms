VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_0rw1r1w_32_512_freepdk45
   CLASS BLOCK ;
   SIZE 237.995 BY 240.69 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  30.5625 0.0 30.7025 0.14 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  33.4225 0.0 33.5625 0.14 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  36.2825 0.0 36.4225 0.14 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  39.1425 0.0 39.2825 0.14 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  42.0025 0.0 42.1425 0.14 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  44.8625 0.0 45.0025 0.14 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  47.7225 0.0 47.8625 0.14 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  50.5825 0.0 50.7225 0.14 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  53.4425 0.0 53.5825 0.14 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  56.3025 0.0 56.4425 0.14 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  59.1625 0.0 59.3025 0.14 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  62.0225 0.0 62.1625 0.14 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  64.8825 0.0 65.0225 0.14 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  67.7425 0.0 67.8825 0.14 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  70.6025 0.0 70.7425 0.14 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  73.4625 0.0 73.6025 0.14 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  76.3225 0.0 76.4625 0.14 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  79.1825 0.0 79.3225 0.14 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  82.0425 0.0 82.1825 0.14 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  84.9025 0.0 85.0425 0.14 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  87.7625 0.0 87.9025 0.14 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  90.6225 0.0 90.7625 0.14 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  93.4825 0.0 93.6225 0.14 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  96.3425 0.0 96.4825 0.14 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  99.2025 0.0 99.3425 0.14 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  102.0625 0.0 102.2025 0.14 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  104.9225 0.0 105.0625 0.14 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  107.7825 0.0 107.9225 0.14 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  110.6425 0.0 110.7825 0.14 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  113.5025 0.0 113.6425 0.14 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  116.3625 0.0 116.5025 0.14 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  119.2225 0.0 119.3625 0.14 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  24.8425 0.0 24.9825 0.14 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  27.7025 0.0 27.8425 0.14 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 57.69 0.14 57.83 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 60.42 0.14 60.56 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 62.63 0.14 62.77 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 65.36 0.14 65.5 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 67.57 0.14 67.71 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 70.3 0.14 70.44 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 72.51 0.14 72.65 ;
      END
   END addr0[8]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  210.1525 240.55 210.2925 240.69 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  207.2925 240.55 207.4325 240.69 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  237.855 25.58 237.995 25.72 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  237.855 22.85 237.995 22.99 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  237.855 20.64 237.995 20.78 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  218.16 0.0 218.3 0.14 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  219.3 0.0 219.44 0.14 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  218.445 0.0 218.585 0.14 ;
      END
   END addr1[7]
   PIN addr1[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  218.73 0.0 218.87 0.14 ;
      END
   END addr1[8]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 7.12 0.14 7.26 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  237.855 234.96 237.995 235.1 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  9.56 0.0 9.7 0.14 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  228.295 240.55 228.435 240.69 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  43.6575 240.55 43.7975 240.69 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  48.3575 240.55 48.4975 240.69 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  53.0575 240.55 53.1975 240.69 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  57.7575 240.55 57.8975 240.69 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  62.4575 240.55 62.5975 240.69 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  67.1575 240.55 67.2975 240.69 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  71.8575 240.55 71.9975 240.69 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  76.5575 240.55 76.6975 240.69 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  81.2575 240.55 81.3975 240.69 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  85.9575 240.55 86.0975 240.69 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  90.6575 240.55 90.7975 240.69 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  95.3575 240.55 95.4975 240.69 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  100.0575 240.55 100.1975 240.69 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  104.7575 240.55 104.8975 240.69 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  109.4575 240.55 109.5975 240.69 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  114.1575 240.55 114.2975 240.69 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  118.8575 240.55 118.9975 240.69 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  123.5575 240.55 123.6975 240.69 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  128.2575 240.55 128.3975 240.69 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  132.9575 240.55 133.0975 240.69 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  137.6575 240.55 137.7975 240.69 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  142.3575 240.55 142.4975 240.69 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  147.0575 240.55 147.1975 240.69 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  151.7575 240.55 151.8975 240.69 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  156.4575 240.55 156.5975 240.69 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  161.1575 240.55 161.2975 240.69 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  165.8575 240.55 165.9975 240.69 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  170.5575 240.55 170.6975 240.69 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  175.2575 240.55 175.3975 240.69 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  179.9575 240.55 180.0975 240.69 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  184.6575 240.55 184.7975 240.69 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  189.3575 240.55 189.4975 240.69 ;
      END
   END dout1[31]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 237.855 240.55 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 237.855 240.55 ;
   LAYER  metal3 ;
      RECT  0.28 57.55 237.855 57.97 ;
      RECT  0.14 57.97 0.28 60.28 ;
      RECT  0.14 60.7 0.28 62.49 ;
      RECT  0.14 62.91 0.28 65.22 ;
      RECT  0.14 65.64 0.28 67.43 ;
      RECT  0.14 67.85 0.28 70.16 ;
      RECT  0.14 70.58 0.28 72.37 ;
      RECT  0.14 72.79 0.28 240.55 ;
      RECT  0.28 0.14 237.715 25.44 ;
      RECT  0.28 25.44 237.715 25.86 ;
      RECT  0.28 25.86 237.715 57.55 ;
      RECT  237.715 25.86 237.855 57.55 ;
      RECT  237.715 23.13 237.855 25.44 ;
      RECT  237.715 0.14 237.855 20.5 ;
      RECT  237.715 20.92 237.855 22.71 ;
      RECT  0.14 0.14 0.28 6.98 ;
      RECT  0.14 7.4 0.28 57.55 ;
      RECT  0.28 57.97 237.715 234.82 ;
      RECT  0.28 234.82 237.715 235.24 ;
      RECT  0.28 235.24 237.715 240.55 ;
      RECT  237.715 57.97 237.855 234.82 ;
      RECT  237.715 235.24 237.855 240.55 ;
   LAYER  metal4 ;
      RECT  0.14 0.42 30.2825 240.55 ;
      RECT  30.2825 0.42 30.9825 240.55 ;
      RECT  30.9825 0.14 33.1425 0.42 ;
      RECT  33.8425 0.14 36.0025 0.42 ;
      RECT  36.7025 0.14 38.8625 0.42 ;
      RECT  39.5625 0.14 41.7225 0.42 ;
      RECT  42.4225 0.14 44.5825 0.42 ;
      RECT  45.2825 0.14 47.4425 0.42 ;
      RECT  48.1425 0.14 50.3025 0.42 ;
      RECT  51.0025 0.14 53.1625 0.42 ;
      RECT  53.8625 0.14 56.0225 0.42 ;
      RECT  56.7225 0.14 58.8825 0.42 ;
      RECT  59.5825 0.14 61.7425 0.42 ;
      RECT  62.4425 0.14 64.6025 0.42 ;
      RECT  65.3025 0.14 67.4625 0.42 ;
      RECT  68.1625 0.14 70.3225 0.42 ;
      RECT  71.0225 0.14 73.1825 0.42 ;
      RECT  73.8825 0.14 76.0425 0.42 ;
      RECT  76.7425 0.14 78.9025 0.42 ;
      RECT  79.6025 0.14 81.7625 0.42 ;
      RECT  82.4625 0.14 84.6225 0.42 ;
      RECT  85.3225 0.14 87.4825 0.42 ;
      RECT  88.1825 0.14 90.3425 0.42 ;
      RECT  91.0425 0.14 93.2025 0.42 ;
      RECT  93.9025 0.14 96.0625 0.42 ;
      RECT  96.7625 0.14 98.9225 0.42 ;
      RECT  99.6225 0.14 101.7825 0.42 ;
      RECT  102.4825 0.14 104.6425 0.42 ;
      RECT  105.3425 0.14 107.5025 0.42 ;
      RECT  108.2025 0.14 110.3625 0.42 ;
      RECT  111.0625 0.14 113.2225 0.42 ;
      RECT  113.9225 0.14 116.0825 0.42 ;
      RECT  116.7825 0.14 118.9425 0.42 ;
      RECT  25.2625 0.14 27.4225 0.42 ;
      RECT  28.1225 0.14 30.2825 0.42 ;
      RECT  30.9825 0.42 209.8725 240.27 ;
      RECT  209.8725 0.42 210.5725 240.27 ;
      RECT  210.5725 0.42 237.855 240.27 ;
      RECT  207.7125 240.27 209.8725 240.55 ;
      RECT  119.6425 0.14 217.88 0.42 ;
      RECT  219.72 0.14 237.855 0.42 ;
      RECT  0.14 0.14 9.28 0.42 ;
      RECT  9.98 0.14 24.5625 0.42 ;
      RECT  210.5725 240.27 228.015 240.55 ;
      RECT  228.715 240.27 237.855 240.55 ;
      RECT  30.9825 240.27 43.3775 240.55 ;
      RECT  44.0775 240.27 48.0775 240.55 ;
      RECT  48.7775 240.27 52.7775 240.55 ;
      RECT  53.4775 240.27 57.4775 240.55 ;
      RECT  58.1775 240.27 62.1775 240.55 ;
      RECT  62.8775 240.27 66.8775 240.55 ;
      RECT  67.5775 240.27 71.5775 240.55 ;
      RECT  72.2775 240.27 76.2775 240.55 ;
      RECT  76.9775 240.27 80.9775 240.55 ;
      RECT  81.6775 240.27 85.6775 240.55 ;
      RECT  86.3775 240.27 90.3775 240.55 ;
      RECT  91.0775 240.27 95.0775 240.55 ;
      RECT  95.7775 240.27 99.7775 240.55 ;
      RECT  100.4775 240.27 104.4775 240.55 ;
      RECT  105.1775 240.27 109.1775 240.55 ;
      RECT  109.8775 240.27 113.8775 240.55 ;
      RECT  114.5775 240.27 118.5775 240.55 ;
      RECT  119.2775 240.27 123.2775 240.55 ;
      RECT  123.9775 240.27 127.9775 240.55 ;
      RECT  128.6775 240.27 132.6775 240.55 ;
      RECT  133.3775 240.27 137.3775 240.55 ;
      RECT  138.0775 240.27 142.0775 240.55 ;
      RECT  142.7775 240.27 146.7775 240.55 ;
      RECT  147.4775 240.27 151.4775 240.55 ;
      RECT  152.1775 240.27 156.1775 240.55 ;
      RECT  156.8775 240.27 160.8775 240.55 ;
      RECT  161.5775 240.27 165.5775 240.55 ;
      RECT  166.2775 240.27 170.2775 240.55 ;
      RECT  170.9775 240.27 174.9775 240.55 ;
      RECT  175.6775 240.27 179.6775 240.55 ;
      RECT  180.3775 240.27 184.3775 240.55 ;
      RECT  185.0775 240.27 189.0775 240.55 ;
      RECT  189.7775 240.27 207.0125 240.55 ;
   END
END    sram_0rw1r1w_32_512_freepdk45
END    LIBRARY
