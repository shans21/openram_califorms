VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_0rw1r1w_512_16_freepdk45
   CLASS BLOCK ;
   SIZE 1589.875 BY 172.25 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  125.7675 0.0 125.9075 0.14 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  128.6275 0.0 128.7675 0.14 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  131.4875 0.0 131.6275 0.14 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  134.3475 0.0 134.4875 0.14 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  137.2075 0.0 137.3475 0.14 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  140.0675 0.0 140.2075 0.14 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  142.9275 0.0 143.0675 0.14 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  145.7875 0.0 145.9275 0.14 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  148.6475 0.0 148.7875 0.14 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  151.5075 0.0 151.6475 0.14 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  154.3675 0.0 154.5075 0.14 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  157.2275 0.0 157.3675 0.14 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  160.0875 0.0 160.2275 0.14 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  162.9475 0.0 163.0875 0.14 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  165.8075 0.0 165.9475 0.14 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  168.6675 0.0 168.8075 0.14 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  171.5275 0.0 171.6675 0.14 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  174.3875 0.0 174.5275 0.14 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  177.2475 0.0 177.3875 0.14 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  180.1075 0.0 180.2475 0.14 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  182.9675 0.0 183.1075 0.14 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  185.8275 0.0 185.9675 0.14 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  188.6875 0.0 188.8275 0.14 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  191.5475 0.0 191.6875 0.14 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  194.4075 0.0 194.5475 0.14 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  197.2675 0.0 197.4075 0.14 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  200.1275 0.0 200.2675 0.14 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  202.9875 0.0 203.1275 0.14 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  205.8475 0.0 205.9875 0.14 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  208.7075 0.0 208.8475 0.14 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  211.5675 0.0 211.7075 0.14 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  214.4275 0.0 214.5675 0.14 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  217.2875 0.0 217.4275 0.14 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  220.1475 0.0 220.2875 0.14 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  223.0075 0.0 223.1475 0.14 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  225.8675 0.0 226.0075 0.14 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  228.7275 0.0 228.8675 0.14 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  231.5875 0.0 231.7275 0.14 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  234.4475 0.0 234.5875 0.14 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  237.3075 0.0 237.4475 0.14 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  240.1675 0.0 240.3075 0.14 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  243.0275 0.0 243.1675 0.14 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  245.8875 0.0 246.0275 0.14 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  248.7475 0.0 248.8875 0.14 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  251.6075 0.0 251.7475 0.14 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  254.4675 0.0 254.6075 0.14 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  257.3275 0.0 257.4675 0.14 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  260.1875 0.0 260.3275 0.14 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  263.0475 0.0 263.1875 0.14 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  265.9075 0.0 266.0475 0.14 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  268.7675 0.0 268.9075 0.14 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  271.6275 0.0 271.7675 0.14 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  274.4875 0.0 274.6275 0.14 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  277.3475 0.0 277.4875 0.14 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  280.2075 0.0 280.3475 0.14 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  283.0675 0.0 283.2075 0.14 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  285.9275 0.0 286.0675 0.14 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  288.7875 0.0 288.9275 0.14 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  291.6475 0.0 291.7875 0.14 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  294.5075 0.0 294.6475 0.14 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  297.3675 0.0 297.5075 0.14 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  300.2275 0.0 300.3675 0.14 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  303.0875 0.0 303.2275 0.14 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  305.9475 0.0 306.0875 0.14 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  308.8075 0.0 308.9475 0.14 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  311.6675 0.0 311.8075 0.14 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  314.5275 0.0 314.6675 0.14 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  317.3875 0.0 317.5275 0.14 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  320.2475 0.0 320.3875 0.14 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  323.1075 0.0 323.2475 0.14 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  325.9675 0.0 326.1075 0.14 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  328.8275 0.0 328.9675 0.14 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  331.6875 0.0 331.8275 0.14 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  334.5475 0.0 334.6875 0.14 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  337.4075 0.0 337.5475 0.14 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  340.2675 0.0 340.4075 0.14 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  343.1275 0.0 343.2675 0.14 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  345.9875 0.0 346.1275 0.14 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  348.8475 0.0 348.9875 0.14 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  351.7075 0.0 351.8475 0.14 ;
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  354.5675 0.0 354.7075 0.14 ;
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  357.4275 0.0 357.5675 0.14 ;
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  360.2875 0.0 360.4275 0.14 ;
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  363.1475 0.0 363.2875 0.14 ;
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  366.0075 0.0 366.1475 0.14 ;
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  368.8675 0.0 369.0075 0.14 ;
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  371.7275 0.0 371.8675 0.14 ;
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  374.5875 0.0 374.7275 0.14 ;
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  377.4475 0.0 377.5875 0.14 ;
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  380.3075 0.0 380.4475 0.14 ;
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  383.1675 0.0 383.3075 0.14 ;
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  386.0275 0.0 386.1675 0.14 ;
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  388.8875 0.0 389.0275 0.14 ;
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  391.7475 0.0 391.8875 0.14 ;
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  394.6075 0.0 394.7475 0.14 ;
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  397.4675 0.0 397.6075 0.14 ;
      END
   END din0[95]
   PIN din0[96]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  400.3275 0.0 400.4675 0.14 ;
      END
   END din0[96]
   PIN din0[97]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  403.1875 0.0 403.3275 0.14 ;
      END
   END din0[97]
   PIN din0[98]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  406.0475 0.0 406.1875 0.14 ;
      END
   END din0[98]
   PIN din0[99]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  408.9075 0.0 409.0475 0.14 ;
      END
   END din0[99]
   PIN din0[100]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  411.7675 0.0 411.9075 0.14 ;
      END
   END din0[100]
   PIN din0[101]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  414.6275 0.0 414.7675 0.14 ;
      END
   END din0[101]
   PIN din0[102]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  417.4875 0.0 417.6275 0.14 ;
      END
   END din0[102]
   PIN din0[103]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  420.3475 0.0 420.4875 0.14 ;
      END
   END din0[103]
   PIN din0[104]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  423.2075 0.0 423.3475 0.14 ;
      END
   END din0[104]
   PIN din0[105]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  426.0675 0.0 426.2075 0.14 ;
      END
   END din0[105]
   PIN din0[106]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  428.9275 0.0 429.0675 0.14 ;
      END
   END din0[106]
   PIN din0[107]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  431.7875 0.0 431.9275 0.14 ;
      END
   END din0[107]
   PIN din0[108]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  434.6475 0.0 434.7875 0.14 ;
      END
   END din0[108]
   PIN din0[109]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  437.5075 0.0 437.6475 0.14 ;
      END
   END din0[109]
   PIN din0[110]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  440.3675 0.0 440.5075 0.14 ;
      END
   END din0[110]
   PIN din0[111]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  443.2275 0.0 443.3675 0.14 ;
      END
   END din0[111]
   PIN din0[112]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  446.0875 0.0 446.2275 0.14 ;
      END
   END din0[112]
   PIN din0[113]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  448.9475 0.0 449.0875 0.14 ;
      END
   END din0[113]
   PIN din0[114]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  451.8075 0.0 451.9475 0.14 ;
      END
   END din0[114]
   PIN din0[115]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  454.6675 0.0 454.8075 0.14 ;
      END
   END din0[115]
   PIN din0[116]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  457.5275 0.0 457.6675 0.14 ;
      END
   END din0[116]
   PIN din0[117]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  460.3875 0.0 460.5275 0.14 ;
      END
   END din0[117]
   PIN din0[118]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  463.2475 0.0 463.3875 0.14 ;
      END
   END din0[118]
   PIN din0[119]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  466.1075 0.0 466.2475 0.14 ;
      END
   END din0[119]
   PIN din0[120]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  468.9675 0.0 469.1075 0.14 ;
      END
   END din0[120]
   PIN din0[121]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  471.8275 0.0 471.9675 0.14 ;
      END
   END din0[121]
   PIN din0[122]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  474.6875 0.0 474.8275 0.14 ;
      END
   END din0[122]
   PIN din0[123]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  477.5475 0.0 477.6875 0.14 ;
      END
   END din0[123]
   PIN din0[124]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  480.4075 0.0 480.5475 0.14 ;
      END
   END din0[124]
   PIN din0[125]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  483.2675 0.0 483.4075 0.14 ;
      END
   END din0[125]
   PIN din0[126]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  486.1275 0.0 486.2675 0.14 ;
      END
   END din0[126]
   PIN din0[127]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  488.9875 0.0 489.1275 0.14 ;
      END
   END din0[127]
   PIN din0[128]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  491.8475 0.0 491.9875 0.14 ;
      END
   END din0[128]
   PIN din0[129]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  494.7075 0.0 494.8475 0.14 ;
      END
   END din0[129]
   PIN din0[130]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  497.5675 0.0 497.7075 0.14 ;
      END
   END din0[130]
   PIN din0[131]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  500.4275 0.0 500.5675 0.14 ;
      END
   END din0[131]
   PIN din0[132]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  503.2875 0.0 503.4275 0.14 ;
      END
   END din0[132]
   PIN din0[133]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  506.1475 0.0 506.2875 0.14 ;
      END
   END din0[133]
   PIN din0[134]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  509.0075 0.0 509.1475 0.14 ;
      END
   END din0[134]
   PIN din0[135]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  511.8675 0.0 512.0075 0.14 ;
      END
   END din0[135]
   PIN din0[136]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  514.7275 0.0 514.8675 0.14 ;
      END
   END din0[136]
   PIN din0[137]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  517.5875 0.0 517.7275 0.14 ;
      END
   END din0[137]
   PIN din0[138]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  520.4475 0.0 520.5875 0.14 ;
      END
   END din0[138]
   PIN din0[139]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  523.3075 0.0 523.4475 0.14 ;
      END
   END din0[139]
   PIN din0[140]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  526.1675 0.0 526.3075 0.14 ;
      END
   END din0[140]
   PIN din0[141]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  529.0275 0.0 529.1675 0.14 ;
      END
   END din0[141]
   PIN din0[142]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  531.8875 0.0 532.0275 0.14 ;
      END
   END din0[142]
   PIN din0[143]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  534.7475 0.0 534.8875 0.14 ;
      END
   END din0[143]
   PIN din0[144]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  537.6075 0.0 537.7475 0.14 ;
      END
   END din0[144]
   PIN din0[145]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  540.4675 0.0 540.6075 0.14 ;
      END
   END din0[145]
   PIN din0[146]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  543.3275 0.0 543.4675 0.14 ;
      END
   END din0[146]
   PIN din0[147]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  546.1875 0.0 546.3275 0.14 ;
      END
   END din0[147]
   PIN din0[148]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  549.0475 0.0 549.1875 0.14 ;
      END
   END din0[148]
   PIN din0[149]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  551.9075 0.0 552.0475 0.14 ;
      END
   END din0[149]
   PIN din0[150]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  554.7675 0.0 554.9075 0.14 ;
      END
   END din0[150]
   PIN din0[151]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  557.6275 0.0 557.7675 0.14 ;
      END
   END din0[151]
   PIN din0[152]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  560.4875 0.0 560.6275 0.14 ;
      END
   END din0[152]
   PIN din0[153]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  563.3475 0.0 563.4875 0.14 ;
      END
   END din0[153]
   PIN din0[154]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  566.2075 0.0 566.3475 0.14 ;
      END
   END din0[154]
   PIN din0[155]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  569.0675 0.0 569.2075 0.14 ;
      END
   END din0[155]
   PIN din0[156]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  571.9275 0.0 572.0675 0.14 ;
      END
   END din0[156]
   PIN din0[157]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  574.7875 0.0 574.9275 0.14 ;
      END
   END din0[157]
   PIN din0[158]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  577.6475 0.0 577.7875 0.14 ;
      END
   END din0[158]
   PIN din0[159]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  580.5075 0.0 580.6475 0.14 ;
      END
   END din0[159]
   PIN din0[160]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  583.3675 0.0 583.5075 0.14 ;
      END
   END din0[160]
   PIN din0[161]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  586.2275 0.0 586.3675 0.14 ;
      END
   END din0[161]
   PIN din0[162]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  589.0875 0.0 589.2275 0.14 ;
      END
   END din0[162]
   PIN din0[163]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  591.9475 0.0 592.0875 0.14 ;
      END
   END din0[163]
   PIN din0[164]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  594.8075 0.0 594.9475 0.14 ;
      END
   END din0[164]
   PIN din0[165]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  597.6675 0.0 597.8075 0.14 ;
      END
   END din0[165]
   PIN din0[166]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  600.5275 0.0 600.6675 0.14 ;
      END
   END din0[166]
   PIN din0[167]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  603.3875 0.0 603.5275 0.14 ;
      END
   END din0[167]
   PIN din0[168]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  606.2475 0.0 606.3875 0.14 ;
      END
   END din0[168]
   PIN din0[169]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  609.1075 0.0 609.2475 0.14 ;
      END
   END din0[169]
   PIN din0[170]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  611.9675 0.0 612.1075 0.14 ;
      END
   END din0[170]
   PIN din0[171]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  614.8275 0.0 614.9675 0.14 ;
      END
   END din0[171]
   PIN din0[172]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  617.6875 0.0 617.8275 0.14 ;
      END
   END din0[172]
   PIN din0[173]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  620.5475 0.0 620.6875 0.14 ;
      END
   END din0[173]
   PIN din0[174]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  623.4075 0.0 623.5475 0.14 ;
      END
   END din0[174]
   PIN din0[175]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  626.2675 0.0 626.4075 0.14 ;
      END
   END din0[175]
   PIN din0[176]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  629.1275 0.0 629.2675 0.14 ;
      END
   END din0[176]
   PIN din0[177]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  631.9875 0.0 632.1275 0.14 ;
      END
   END din0[177]
   PIN din0[178]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  634.8475 0.0 634.9875 0.14 ;
      END
   END din0[178]
   PIN din0[179]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  637.7075 0.0 637.8475 0.14 ;
      END
   END din0[179]
   PIN din0[180]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  640.5675 0.0 640.7075 0.14 ;
      END
   END din0[180]
   PIN din0[181]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  643.4275 0.0 643.5675 0.14 ;
      END
   END din0[181]
   PIN din0[182]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  646.2875 0.0 646.4275 0.14 ;
      END
   END din0[182]
   PIN din0[183]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  649.1475 0.0 649.2875 0.14 ;
      END
   END din0[183]
   PIN din0[184]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  652.0075 0.0 652.1475 0.14 ;
      END
   END din0[184]
   PIN din0[185]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  654.8675 0.0 655.0075 0.14 ;
      END
   END din0[185]
   PIN din0[186]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  657.7275 0.0 657.8675 0.14 ;
      END
   END din0[186]
   PIN din0[187]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  660.5875 0.0 660.7275 0.14 ;
      END
   END din0[187]
   PIN din0[188]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  663.4475 0.0 663.5875 0.14 ;
      END
   END din0[188]
   PIN din0[189]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  666.3075 0.0 666.4475 0.14 ;
      END
   END din0[189]
   PIN din0[190]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  669.1675 0.0 669.3075 0.14 ;
      END
   END din0[190]
   PIN din0[191]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  672.0275 0.0 672.1675 0.14 ;
      END
   END din0[191]
   PIN din0[192]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  674.8875 0.0 675.0275 0.14 ;
      END
   END din0[192]
   PIN din0[193]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  677.7475 0.0 677.8875 0.14 ;
      END
   END din0[193]
   PIN din0[194]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  680.6075 0.0 680.7475 0.14 ;
      END
   END din0[194]
   PIN din0[195]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  683.4675 0.0 683.6075 0.14 ;
      END
   END din0[195]
   PIN din0[196]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  686.3275 0.0 686.4675 0.14 ;
      END
   END din0[196]
   PIN din0[197]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  689.1875 0.0 689.3275 0.14 ;
      END
   END din0[197]
   PIN din0[198]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  692.0475 0.0 692.1875 0.14 ;
      END
   END din0[198]
   PIN din0[199]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  694.9075 0.0 695.0475 0.14 ;
      END
   END din0[199]
   PIN din0[200]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  697.7675 0.0 697.9075 0.14 ;
      END
   END din0[200]
   PIN din0[201]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  700.6275 0.0 700.7675 0.14 ;
      END
   END din0[201]
   PIN din0[202]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  703.4875 0.0 703.6275 0.14 ;
      END
   END din0[202]
   PIN din0[203]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  706.3475 0.0 706.4875 0.14 ;
      END
   END din0[203]
   PIN din0[204]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  709.2075 0.0 709.3475 0.14 ;
      END
   END din0[204]
   PIN din0[205]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  712.0675 0.0 712.2075 0.14 ;
      END
   END din0[205]
   PIN din0[206]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  714.9275 0.0 715.0675 0.14 ;
      END
   END din0[206]
   PIN din0[207]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  717.7875 0.0 717.9275 0.14 ;
      END
   END din0[207]
   PIN din0[208]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  720.6475 0.0 720.7875 0.14 ;
      END
   END din0[208]
   PIN din0[209]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  723.5075 0.0 723.6475 0.14 ;
      END
   END din0[209]
   PIN din0[210]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  726.3675 0.0 726.5075 0.14 ;
      END
   END din0[210]
   PIN din0[211]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  729.2275 0.0 729.3675 0.14 ;
      END
   END din0[211]
   PIN din0[212]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  732.0875 0.0 732.2275 0.14 ;
      END
   END din0[212]
   PIN din0[213]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  734.9475 0.0 735.0875 0.14 ;
      END
   END din0[213]
   PIN din0[214]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  737.8075 0.0 737.9475 0.14 ;
      END
   END din0[214]
   PIN din0[215]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  740.6675 0.0 740.8075 0.14 ;
      END
   END din0[215]
   PIN din0[216]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  743.5275 0.0 743.6675 0.14 ;
      END
   END din0[216]
   PIN din0[217]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  746.3875 0.0 746.5275 0.14 ;
      END
   END din0[217]
   PIN din0[218]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  749.2475 0.0 749.3875 0.14 ;
      END
   END din0[218]
   PIN din0[219]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  752.1075 0.0 752.2475 0.14 ;
      END
   END din0[219]
   PIN din0[220]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  754.9675 0.0 755.1075 0.14 ;
      END
   END din0[220]
   PIN din0[221]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  757.8275 0.0 757.9675 0.14 ;
      END
   END din0[221]
   PIN din0[222]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  760.6875 0.0 760.8275 0.14 ;
      END
   END din0[222]
   PIN din0[223]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  763.5475 0.0 763.6875 0.14 ;
      END
   END din0[223]
   PIN din0[224]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  766.4075 0.0 766.5475 0.14 ;
      END
   END din0[224]
   PIN din0[225]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  769.2675 0.0 769.4075 0.14 ;
      END
   END din0[225]
   PIN din0[226]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  772.1275 0.0 772.2675 0.14 ;
      END
   END din0[226]
   PIN din0[227]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  774.9875 0.0 775.1275 0.14 ;
      END
   END din0[227]
   PIN din0[228]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  777.8475 0.0 777.9875 0.14 ;
      END
   END din0[228]
   PIN din0[229]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  780.7075 0.0 780.8475 0.14 ;
      END
   END din0[229]
   PIN din0[230]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  783.5675 0.0 783.7075 0.14 ;
      END
   END din0[230]
   PIN din0[231]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  786.4275 0.0 786.5675 0.14 ;
      END
   END din0[231]
   PIN din0[232]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  789.2875 0.0 789.4275 0.14 ;
      END
   END din0[232]
   PIN din0[233]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  792.1475 0.0 792.2875 0.14 ;
      END
   END din0[233]
   PIN din0[234]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  795.0075 0.0 795.1475 0.14 ;
      END
   END din0[234]
   PIN din0[235]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  797.8675 0.0 798.0075 0.14 ;
      END
   END din0[235]
   PIN din0[236]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  800.7275 0.0 800.8675 0.14 ;
      END
   END din0[236]
   PIN din0[237]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  803.5875 0.0 803.7275 0.14 ;
      END
   END din0[237]
   PIN din0[238]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  806.4475 0.0 806.5875 0.14 ;
      END
   END din0[238]
   PIN din0[239]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  809.3075 0.0 809.4475 0.14 ;
      END
   END din0[239]
   PIN din0[240]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  812.1675 0.0 812.3075 0.14 ;
      END
   END din0[240]
   PIN din0[241]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  815.0275 0.0 815.1675 0.14 ;
      END
   END din0[241]
   PIN din0[242]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  817.8875 0.0 818.0275 0.14 ;
      END
   END din0[242]
   PIN din0[243]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  820.7475 0.0 820.8875 0.14 ;
      END
   END din0[243]
   PIN din0[244]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  823.6075 0.0 823.7475 0.14 ;
      END
   END din0[244]
   PIN din0[245]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  826.4675 0.0 826.6075 0.14 ;
      END
   END din0[245]
   PIN din0[246]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  829.3275 0.0 829.4675 0.14 ;
      END
   END din0[246]
   PIN din0[247]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  832.1875 0.0 832.3275 0.14 ;
      END
   END din0[247]
   PIN din0[248]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  835.0475 0.0 835.1875 0.14 ;
      END
   END din0[248]
   PIN din0[249]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  837.9075 0.0 838.0475 0.14 ;
      END
   END din0[249]
   PIN din0[250]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  840.7675 0.0 840.9075 0.14 ;
      END
   END din0[250]
   PIN din0[251]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  843.6275 0.0 843.7675 0.14 ;
      END
   END din0[251]
   PIN din0[252]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  846.4875 0.0 846.6275 0.14 ;
      END
   END din0[252]
   PIN din0[253]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  849.3475 0.0 849.4875 0.14 ;
      END
   END din0[253]
   PIN din0[254]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  852.2075 0.0 852.3475 0.14 ;
      END
   END din0[254]
   PIN din0[255]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  855.0675 0.0 855.2075 0.14 ;
      END
   END din0[255]
   PIN din0[256]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  857.9275 0.0 858.0675 0.14 ;
      END
   END din0[256]
   PIN din0[257]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  860.7875 0.0 860.9275 0.14 ;
      END
   END din0[257]
   PIN din0[258]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  863.6475 0.0 863.7875 0.14 ;
      END
   END din0[258]
   PIN din0[259]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  866.5075 0.0 866.6475 0.14 ;
      END
   END din0[259]
   PIN din0[260]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  869.3675 0.0 869.5075 0.14 ;
      END
   END din0[260]
   PIN din0[261]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  872.2275 0.0 872.3675 0.14 ;
      END
   END din0[261]
   PIN din0[262]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  875.0875 0.0 875.2275 0.14 ;
      END
   END din0[262]
   PIN din0[263]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  877.9475 0.0 878.0875 0.14 ;
      END
   END din0[263]
   PIN din0[264]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  880.8075 0.0 880.9475 0.14 ;
      END
   END din0[264]
   PIN din0[265]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  883.6675 0.0 883.8075 0.14 ;
      END
   END din0[265]
   PIN din0[266]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  886.5275 0.0 886.6675 0.14 ;
      END
   END din0[266]
   PIN din0[267]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  889.3875 0.0 889.5275 0.14 ;
      END
   END din0[267]
   PIN din0[268]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  892.2475 0.0 892.3875 0.14 ;
      END
   END din0[268]
   PIN din0[269]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  895.1075 0.0 895.2475 0.14 ;
      END
   END din0[269]
   PIN din0[270]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  897.9675 0.0 898.1075 0.14 ;
      END
   END din0[270]
   PIN din0[271]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  900.8275 0.0 900.9675 0.14 ;
      END
   END din0[271]
   PIN din0[272]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  903.6875 0.0 903.8275 0.14 ;
      END
   END din0[272]
   PIN din0[273]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  906.5475 0.0 906.6875 0.14 ;
      END
   END din0[273]
   PIN din0[274]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  909.4075 0.0 909.5475 0.14 ;
      END
   END din0[274]
   PIN din0[275]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  912.2675 0.0 912.4075 0.14 ;
      END
   END din0[275]
   PIN din0[276]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  915.1275 0.0 915.2675 0.14 ;
      END
   END din0[276]
   PIN din0[277]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  917.9875 0.0 918.1275 0.14 ;
      END
   END din0[277]
   PIN din0[278]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  920.8475 0.0 920.9875 0.14 ;
      END
   END din0[278]
   PIN din0[279]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  923.7075 0.0 923.8475 0.14 ;
      END
   END din0[279]
   PIN din0[280]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  926.5675 0.0 926.7075 0.14 ;
      END
   END din0[280]
   PIN din0[281]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  929.4275 0.0 929.5675 0.14 ;
      END
   END din0[281]
   PIN din0[282]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  932.2875 0.0 932.4275 0.14 ;
      END
   END din0[282]
   PIN din0[283]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  935.1475 0.0 935.2875 0.14 ;
      END
   END din0[283]
   PIN din0[284]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  938.0075 0.0 938.1475 0.14 ;
      END
   END din0[284]
   PIN din0[285]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  940.8675 0.0 941.0075 0.14 ;
      END
   END din0[285]
   PIN din0[286]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  943.7275 0.0 943.8675 0.14 ;
      END
   END din0[286]
   PIN din0[287]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  946.5875 0.0 946.7275 0.14 ;
      END
   END din0[287]
   PIN din0[288]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  949.4475 0.0 949.5875 0.14 ;
      END
   END din0[288]
   PIN din0[289]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  952.3075 0.0 952.4475 0.14 ;
      END
   END din0[289]
   PIN din0[290]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  955.1675 0.0 955.3075 0.14 ;
      END
   END din0[290]
   PIN din0[291]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  958.0275 0.0 958.1675 0.14 ;
      END
   END din0[291]
   PIN din0[292]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  960.8875 0.0 961.0275 0.14 ;
      END
   END din0[292]
   PIN din0[293]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  963.7475 0.0 963.8875 0.14 ;
      END
   END din0[293]
   PIN din0[294]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  966.6075 0.0 966.7475 0.14 ;
      END
   END din0[294]
   PIN din0[295]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  969.4675 0.0 969.6075 0.14 ;
      END
   END din0[295]
   PIN din0[296]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  972.3275 0.0 972.4675 0.14 ;
      END
   END din0[296]
   PIN din0[297]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  975.1875 0.0 975.3275 0.14 ;
      END
   END din0[297]
   PIN din0[298]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  978.0475 0.0 978.1875 0.14 ;
      END
   END din0[298]
   PIN din0[299]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  980.9075 0.0 981.0475 0.14 ;
      END
   END din0[299]
   PIN din0[300]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  983.7675 0.0 983.9075 0.14 ;
      END
   END din0[300]
   PIN din0[301]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  986.6275 0.0 986.7675 0.14 ;
      END
   END din0[301]
   PIN din0[302]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  989.4875 0.0 989.6275 0.14 ;
      END
   END din0[302]
   PIN din0[303]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  992.3475 0.0 992.4875 0.14 ;
      END
   END din0[303]
   PIN din0[304]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  995.2075 0.0 995.3475 0.14 ;
      END
   END din0[304]
   PIN din0[305]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  998.0675 0.0 998.2075 0.14 ;
      END
   END din0[305]
   PIN din0[306]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1000.9275 0.0 1001.0675 0.14 ;
      END
   END din0[306]
   PIN din0[307]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1003.7875 0.0 1003.9275 0.14 ;
      END
   END din0[307]
   PIN din0[308]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1006.6475 0.0 1006.7875 0.14 ;
      END
   END din0[308]
   PIN din0[309]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1009.5075 0.0 1009.6475 0.14 ;
      END
   END din0[309]
   PIN din0[310]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1012.3675 0.0 1012.5075 0.14 ;
      END
   END din0[310]
   PIN din0[311]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1015.2275 0.0 1015.3675 0.14 ;
      END
   END din0[311]
   PIN din0[312]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1018.0875 0.0 1018.2275 0.14 ;
      END
   END din0[312]
   PIN din0[313]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1020.9475 0.0 1021.0875 0.14 ;
      END
   END din0[313]
   PIN din0[314]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1023.8075 0.0 1023.9475 0.14 ;
      END
   END din0[314]
   PIN din0[315]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1026.6675 0.0 1026.8075 0.14 ;
      END
   END din0[315]
   PIN din0[316]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1029.5275 0.0 1029.6675 0.14 ;
      END
   END din0[316]
   PIN din0[317]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1032.3875 0.0 1032.5275 0.14 ;
      END
   END din0[317]
   PIN din0[318]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1035.2475 0.0 1035.3875 0.14 ;
      END
   END din0[318]
   PIN din0[319]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1038.1075 0.0 1038.2475 0.14 ;
      END
   END din0[319]
   PIN din0[320]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1040.9675 0.0 1041.1075 0.14 ;
      END
   END din0[320]
   PIN din0[321]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1043.8275 0.0 1043.9675 0.14 ;
      END
   END din0[321]
   PIN din0[322]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1046.6875 0.0 1046.8275 0.14 ;
      END
   END din0[322]
   PIN din0[323]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1049.5475 0.0 1049.6875 0.14 ;
      END
   END din0[323]
   PIN din0[324]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1052.4075 0.0 1052.5475 0.14 ;
      END
   END din0[324]
   PIN din0[325]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1055.2675 0.0 1055.4075 0.14 ;
      END
   END din0[325]
   PIN din0[326]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1058.1275 0.0 1058.2675 0.14 ;
      END
   END din0[326]
   PIN din0[327]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1060.9875 0.0 1061.1275 0.14 ;
      END
   END din0[327]
   PIN din0[328]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1063.8475 0.0 1063.9875 0.14 ;
      END
   END din0[328]
   PIN din0[329]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1066.7075 0.0 1066.8475 0.14 ;
      END
   END din0[329]
   PIN din0[330]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1069.5675 0.0 1069.7075 0.14 ;
      END
   END din0[330]
   PIN din0[331]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1072.4275 0.0 1072.5675 0.14 ;
      END
   END din0[331]
   PIN din0[332]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1075.2875 0.0 1075.4275 0.14 ;
      END
   END din0[332]
   PIN din0[333]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1078.1475 0.0 1078.2875 0.14 ;
      END
   END din0[333]
   PIN din0[334]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1081.0075 0.0 1081.1475 0.14 ;
      END
   END din0[334]
   PIN din0[335]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1083.8675 0.0 1084.0075 0.14 ;
      END
   END din0[335]
   PIN din0[336]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1086.7275 0.0 1086.8675 0.14 ;
      END
   END din0[336]
   PIN din0[337]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1089.5875 0.0 1089.7275 0.14 ;
      END
   END din0[337]
   PIN din0[338]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1092.4475 0.0 1092.5875 0.14 ;
      END
   END din0[338]
   PIN din0[339]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1095.3075 0.0 1095.4475 0.14 ;
      END
   END din0[339]
   PIN din0[340]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1098.1675 0.0 1098.3075 0.14 ;
      END
   END din0[340]
   PIN din0[341]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1101.0275 0.0 1101.1675 0.14 ;
      END
   END din0[341]
   PIN din0[342]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1103.8875 0.0 1104.0275 0.14 ;
      END
   END din0[342]
   PIN din0[343]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1106.7475 0.0 1106.8875 0.14 ;
      END
   END din0[343]
   PIN din0[344]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1109.6075 0.0 1109.7475 0.14 ;
      END
   END din0[344]
   PIN din0[345]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1112.4675 0.0 1112.6075 0.14 ;
      END
   END din0[345]
   PIN din0[346]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1115.3275 0.0 1115.4675 0.14 ;
      END
   END din0[346]
   PIN din0[347]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1118.1875 0.0 1118.3275 0.14 ;
      END
   END din0[347]
   PIN din0[348]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1121.0475 0.0 1121.1875 0.14 ;
      END
   END din0[348]
   PIN din0[349]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1123.9075 0.0 1124.0475 0.14 ;
      END
   END din0[349]
   PIN din0[350]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1126.7675 0.0 1126.9075 0.14 ;
      END
   END din0[350]
   PIN din0[351]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1129.6275 0.0 1129.7675 0.14 ;
      END
   END din0[351]
   PIN din0[352]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1132.4875 0.0 1132.6275 0.14 ;
      END
   END din0[352]
   PIN din0[353]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1135.3475 0.0 1135.4875 0.14 ;
      END
   END din0[353]
   PIN din0[354]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1138.2075 0.0 1138.3475 0.14 ;
      END
   END din0[354]
   PIN din0[355]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1141.0675 0.0 1141.2075 0.14 ;
      END
   END din0[355]
   PIN din0[356]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1143.9275 0.0 1144.0675 0.14 ;
      END
   END din0[356]
   PIN din0[357]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1146.7875 0.0 1146.9275 0.14 ;
      END
   END din0[357]
   PIN din0[358]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1149.6475 0.0 1149.7875 0.14 ;
      END
   END din0[358]
   PIN din0[359]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1152.5075 0.0 1152.6475 0.14 ;
      END
   END din0[359]
   PIN din0[360]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1155.3675 0.0 1155.5075 0.14 ;
      END
   END din0[360]
   PIN din0[361]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1158.2275 0.0 1158.3675 0.14 ;
      END
   END din0[361]
   PIN din0[362]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1161.0875 0.0 1161.2275 0.14 ;
      END
   END din0[362]
   PIN din0[363]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1163.9475 0.0 1164.0875 0.14 ;
      END
   END din0[363]
   PIN din0[364]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1166.8075 0.0 1166.9475 0.14 ;
      END
   END din0[364]
   PIN din0[365]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1169.6675 0.0 1169.8075 0.14 ;
      END
   END din0[365]
   PIN din0[366]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1172.5275 0.0 1172.6675 0.14 ;
      END
   END din0[366]
   PIN din0[367]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1175.3875 0.0 1175.5275 0.14 ;
      END
   END din0[367]
   PIN din0[368]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1178.2475 0.0 1178.3875 0.14 ;
      END
   END din0[368]
   PIN din0[369]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1181.1075 0.0 1181.2475 0.14 ;
      END
   END din0[369]
   PIN din0[370]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1183.9675 0.0 1184.1075 0.14 ;
      END
   END din0[370]
   PIN din0[371]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1186.8275 0.0 1186.9675 0.14 ;
      END
   END din0[371]
   PIN din0[372]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1189.6875 0.0 1189.8275 0.14 ;
      END
   END din0[372]
   PIN din0[373]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1192.5475 0.0 1192.6875 0.14 ;
      END
   END din0[373]
   PIN din0[374]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1195.4075 0.0 1195.5475 0.14 ;
      END
   END din0[374]
   PIN din0[375]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1198.2675 0.0 1198.4075 0.14 ;
      END
   END din0[375]
   PIN din0[376]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1201.1275 0.0 1201.2675 0.14 ;
      END
   END din0[376]
   PIN din0[377]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1203.9875 0.0 1204.1275 0.14 ;
      END
   END din0[377]
   PIN din0[378]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1206.8475 0.0 1206.9875 0.14 ;
      END
   END din0[378]
   PIN din0[379]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1209.7075 0.0 1209.8475 0.14 ;
      END
   END din0[379]
   PIN din0[380]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1212.5675 0.0 1212.7075 0.14 ;
      END
   END din0[380]
   PIN din0[381]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1215.4275 0.0 1215.5675 0.14 ;
      END
   END din0[381]
   PIN din0[382]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1218.2875 0.0 1218.4275 0.14 ;
      END
   END din0[382]
   PIN din0[383]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1221.1475 0.0 1221.2875 0.14 ;
      END
   END din0[383]
   PIN din0[384]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1224.0075 0.0 1224.1475 0.14 ;
      END
   END din0[384]
   PIN din0[385]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1226.8675 0.0 1227.0075 0.14 ;
      END
   END din0[385]
   PIN din0[386]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1229.7275 0.0 1229.8675 0.14 ;
      END
   END din0[386]
   PIN din0[387]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1232.5875 0.0 1232.7275 0.14 ;
      END
   END din0[387]
   PIN din0[388]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1235.4475 0.0 1235.5875 0.14 ;
      END
   END din0[388]
   PIN din0[389]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1238.3075 0.0 1238.4475 0.14 ;
      END
   END din0[389]
   PIN din0[390]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1241.1675 0.0 1241.3075 0.14 ;
      END
   END din0[390]
   PIN din0[391]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1244.0275 0.0 1244.1675 0.14 ;
      END
   END din0[391]
   PIN din0[392]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1246.8875 0.0 1247.0275 0.14 ;
      END
   END din0[392]
   PIN din0[393]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1249.7475 0.0 1249.8875 0.14 ;
      END
   END din0[393]
   PIN din0[394]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1252.6075 0.0 1252.7475 0.14 ;
      END
   END din0[394]
   PIN din0[395]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1255.4675 0.0 1255.6075 0.14 ;
      END
   END din0[395]
   PIN din0[396]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1258.3275 0.0 1258.4675 0.14 ;
      END
   END din0[396]
   PIN din0[397]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1261.1875 0.0 1261.3275 0.14 ;
      END
   END din0[397]
   PIN din0[398]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1264.0475 0.0 1264.1875 0.14 ;
      END
   END din0[398]
   PIN din0[399]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1266.9075 0.0 1267.0475 0.14 ;
      END
   END din0[399]
   PIN din0[400]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1269.7675 0.0 1269.9075 0.14 ;
      END
   END din0[400]
   PIN din0[401]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1272.6275 0.0 1272.7675 0.14 ;
      END
   END din0[401]
   PIN din0[402]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1275.4875 0.0 1275.6275 0.14 ;
      END
   END din0[402]
   PIN din0[403]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1278.3475 0.0 1278.4875 0.14 ;
      END
   END din0[403]
   PIN din0[404]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1281.2075 0.0 1281.3475 0.14 ;
      END
   END din0[404]
   PIN din0[405]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1284.0675 0.0 1284.2075 0.14 ;
      END
   END din0[405]
   PIN din0[406]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1286.9275 0.0 1287.0675 0.14 ;
      END
   END din0[406]
   PIN din0[407]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1289.7875 0.0 1289.9275 0.14 ;
      END
   END din0[407]
   PIN din0[408]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1292.6475 0.0 1292.7875 0.14 ;
      END
   END din0[408]
   PIN din0[409]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1295.5075 0.0 1295.6475 0.14 ;
      END
   END din0[409]
   PIN din0[410]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1298.3675 0.0 1298.5075 0.14 ;
      END
   END din0[410]
   PIN din0[411]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1301.2275 0.0 1301.3675 0.14 ;
      END
   END din0[411]
   PIN din0[412]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1304.0875 0.0 1304.2275 0.14 ;
      END
   END din0[412]
   PIN din0[413]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1306.9475 0.0 1307.0875 0.14 ;
      END
   END din0[413]
   PIN din0[414]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1309.8075 0.0 1309.9475 0.14 ;
      END
   END din0[414]
   PIN din0[415]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1312.6675 0.0 1312.8075 0.14 ;
      END
   END din0[415]
   PIN din0[416]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1315.5275 0.0 1315.6675 0.14 ;
      END
   END din0[416]
   PIN din0[417]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1318.3875 0.0 1318.5275 0.14 ;
      END
   END din0[417]
   PIN din0[418]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1321.2475 0.0 1321.3875 0.14 ;
      END
   END din0[418]
   PIN din0[419]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1324.1075 0.0 1324.2475 0.14 ;
      END
   END din0[419]
   PIN din0[420]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1326.9675 0.0 1327.1075 0.14 ;
      END
   END din0[420]
   PIN din0[421]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1329.8275 0.0 1329.9675 0.14 ;
      END
   END din0[421]
   PIN din0[422]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1332.6875 0.0 1332.8275 0.14 ;
      END
   END din0[422]
   PIN din0[423]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1335.5475 0.0 1335.6875 0.14 ;
      END
   END din0[423]
   PIN din0[424]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1338.4075 0.0 1338.5475 0.14 ;
      END
   END din0[424]
   PIN din0[425]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1341.2675 0.0 1341.4075 0.14 ;
      END
   END din0[425]
   PIN din0[426]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1344.1275 0.0 1344.2675 0.14 ;
      END
   END din0[426]
   PIN din0[427]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1346.9875 0.0 1347.1275 0.14 ;
      END
   END din0[427]
   PIN din0[428]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1349.8475 0.0 1349.9875 0.14 ;
      END
   END din0[428]
   PIN din0[429]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1352.7075 0.0 1352.8475 0.14 ;
      END
   END din0[429]
   PIN din0[430]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1355.5675 0.0 1355.7075 0.14 ;
      END
   END din0[430]
   PIN din0[431]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1358.4275 0.0 1358.5675 0.14 ;
      END
   END din0[431]
   PIN din0[432]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1361.2875 0.0 1361.4275 0.14 ;
      END
   END din0[432]
   PIN din0[433]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1364.1475 0.0 1364.2875 0.14 ;
      END
   END din0[433]
   PIN din0[434]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1367.0075 0.0 1367.1475 0.14 ;
      END
   END din0[434]
   PIN din0[435]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1369.8675 0.0 1370.0075 0.14 ;
      END
   END din0[435]
   PIN din0[436]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1372.7275 0.0 1372.8675 0.14 ;
      END
   END din0[436]
   PIN din0[437]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1375.5875 0.0 1375.7275 0.14 ;
      END
   END din0[437]
   PIN din0[438]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1378.4475 0.0 1378.5875 0.14 ;
      END
   END din0[438]
   PIN din0[439]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1381.3075 0.0 1381.4475 0.14 ;
      END
   END din0[439]
   PIN din0[440]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1384.1675 0.0 1384.3075 0.14 ;
      END
   END din0[440]
   PIN din0[441]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1387.0275 0.0 1387.1675 0.14 ;
      END
   END din0[441]
   PIN din0[442]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1389.8875 0.0 1390.0275 0.14 ;
      END
   END din0[442]
   PIN din0[443]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1392.7475 0.0 1392.8875 0.14 ;
      END
   END din0[443]
   PIN din0[444]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1395.6075 0.0 1395.7475 0.14 ;
      END
   END din0[444]
   PIN din0[445]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1398.4675 0.0 1398.6075 0.14 ;
      END
   END din0[445]
   PIN din0[446]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1401.3275 0.0 1401.4675 0.14 ;
      END
   END din0[446]
   PIN din0[447]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1404.1875 0.0 1404.3275 0.14 ;
      END
   END din0[447]
   PIN din0[448]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1407.0475 0.0 1407.1875 0.14 ;
      END
   END din0[448]
   PIN din0[449]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1409.9075 0.0 1410.0475 0.14 ;
      END
   END din0[449]
   PIN din0[450]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1412.7675 0.0 1412.9075 0.14 ;
      END
   END din0[450]
   PIN din0[451]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1415.6275 0.0 1415.7675 0.14 ;
      END
   END din0[451]
   PIN din0[452]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1418.4875 0.0 1418.6275 0.14 ;
      END
   END din0[452]
   PIN din0[453]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1421.3475 0.0 1421.4875 0.14 ;
      END
   END din0[453]
   PIN din0[454]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1424.2075 0.0 1424.3475 0.14 ;
      END
   END din0[454]
   PIN din0[455]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1427.0675 0.0 1427.2075 0.14 ;
      END
   END din0[455]
   PIN din0[456]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1429.9275 0.0 1430.0675 0.14 ;
      END
   END din0[456]
   PIN din0[457]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1432.7875 0.0 1432.9275 0.14 ;
      END
   END din0[457]
   PIN din0[458]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1435.6475 0.0 1435.7875 0.14 ;
      END
   END din0[458]
   PIN din0[459]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1438.5075 0.0 1438.6475 0.14 ;
      END
   END din0[459]
   PIN din0[460]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1441.3675 0.0 1441.5075 0.14 ;
      END
   END din0[460]
   PIN din0[461]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1444.2275 0.0 1444.3675 0.14 ;
      END
   END din0[461]
   PIN din0[462]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1447.0875 0.0 1447.2275 0.14 ;
      END
   END din0[462]
   PIN din0[463]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1449.9475 0.0 1450.0875 0.14 ;
      END
   END din0[463]
   PIN din0[464]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1452.8075 0.0 1452.9475 0.14 ;
      END
   END din0[464]
   PIN din0[465]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1455.6675 0.0 1455.8075 0.14 ;
      END
   END din0[465]
   PIN din0[466]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1458.5275 0.0 1458.6675 0.14 ;
      END
   END din0[466]
   PIN din0[467]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1461.3875 0.0 1461.5275 0.14 ;
      END
   END din0[467]
   PIN din0[468]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1464.2475 0.0 1464.3875 0.14 ;
      END
   END din0[468]
   PIN din0[469]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1467.1075 0.0 1467.2475 0.14 ;
      END
   END din0[469]
   PIN din0[470]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1469.9675 0.0 1470.1075 0.14 ;
      END
   END din0[470]
   PIN din0[471]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1472.8275 0.0 1472.9675 0.14 ;
      END
   END din0[471]
   PIN din0[472]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1475.6875 0.0 1475.8275 0.14 ;
      END
   END din0[472]
   PIN din0[473]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1478.5475 0.0 1478.6875 0.14 ;
      END
   END din0[473]
   PIN din0[474]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1481.4075 0.0 1481.5475 0.14 ;
      END
   END din0[474]
   PIN din0[475]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1484.2675 0.0 1484.4075 0.14 ;
      END
   END din0[475]
   PIN din0[476]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1487.1275 0.0 1487.2675 0.14 ;
      END
   END din0[476]
   PIN din0[477]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1489.9875 0.0 1490.1275 0.14 ;
      END
   END din0[477]
   PIN din0[478]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1492.8475 0.0 1492.9875 0.14 ;
      END
   END din0[478]
   PIN din0[479]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1495.7075 0.0 1495.8475 0.14 ;
      END
   END din0[479]
   PIN din0[480]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1498.5675 0.0 1498.7075 0.14 ;
      END
   END din0[480]
   PIN din0[481]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1501.4275 0.0 1501.5675 0.14 ;
      END
   END din0[481]
   PIN din0[482]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1504.2875 0.0 1504.4275 0.14 ;
      END
   END din0[482]
   PIN din0[483]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1507.1475 0.0 1507.2875 0.14 ;
      END
   END din0[483]
   PIN din0[484]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1510.0075 0.0 1510.1475 0.14 ;
      END
   END din0[484]
   PIN din0[485]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1512.8675 0.0 1513.0075 0.14 ;
      END
   END din0[485]
   PIN din0[486]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1515.7275 0.0 1515.8675 0.14 ;
      END
   END din0[486]
   PIN din0[487]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1518.5875 0.0 1518.7275 0.14 ;
      END
   END din0[487]
   PIN din0[488]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1521.4475 0.0 1521.5875 0.14 ;
      END
   END din0[488]
   PIN din0[489]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1524.3075 0.0 1524.4475 0.14 ;
      END
   END din0[489]
   PIN din0[490]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1527.1675 0.0 1527.3075 0.14 ;
      END
   END din0[490]
   PIN din0[491]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1530.0275 0.0 1530.1675 0.14 ;
      END
   END din0[491]
   PIN din0[492]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1532.8875 0.0 1533.0275 0.14 ;
      END
   END din0[492]
   PIN din0[493]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1535.7475 0.0 1535.8875 0.14 ;
      END
   END din0[493]
   PIN din0[494]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1538.6075 0.0 1538.7475 0.14 ;
      END
   END din0[494]
   PIN din0[495]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1541.4675 0.0 1541.6075 0.14 ;
      END
   END din0[495]
   PIN din0[496]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1544.3275 0.0 1544.4675 0.14 ;
      END
   END din0[496]
   PIN din0[497]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1547.1875 0.0 1547.3275 0.14 ;
      END
   END din0[497]
   PIN din0[498]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1550.0475 0.0 1550.1875 0.14 ;
      END
   END din0[498]
   PIN din0[499]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1552.9075 0.0 1553.0475 0.14 ;
      END
   END din0[499]
   PIN din0[500]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1555.7675 0.0 1555.9075 0.14 ;
      END
   END din0[500]
   PIN din0[501]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1558.6275 0.0 1558.7675 0.14 ;
      END
   END din0[501]
   PIN din0[502]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1561.4875 0.0 1561.6275 0.14 ;
      END
   END din0[502]
   PIN din0[503]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1564.3475 0.0 1564.4875 0.14 ;
      END
   END din0[503]
   PIN din0[504]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1567.2075 0.0 1567.3475 0.14 ;
      END
   END din0[504]
   PIN din0[505]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1570.0675 0.0 1570.2075 0.14 ;
      END
   END din0[505]
   PIN din0[506]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1572.9275 0.0 1573.0675 0.14 ;
      END
   END din0[506]
   PIN din0[507]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1575.7875 0.0 1575.9275 0.14 ;
      END
   END din0[507]
   PIN din0[508]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1578.6475 0.0 1578.7875 0.14 ;
      END
   END din0[508]
   PIN din0[509]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1581.5075 0.0 1581.6475 0.14 ;
      END
   END din0[509]
   PIN din0[510]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1584.3675 0.0 1584.5075 0.14 ;
      END
   END din0[510]
   PIN din0[511]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1587.2275 0.0 1587.3675 0.14 ;
      END
   END din0[511]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  120.62 172.11 120.76 172.25 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  119.48 172.11 119.62 172.25 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  120.335 172.11 120.475 172.25 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  120.05 172.11 120.19 172.25 ;
      END
   END addr0[3]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  798.555 172.11 798.695 172.25 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  798.27 172.11 798.41 172.25 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  799.125 172.11 799.265 172.25 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  798.5575 172.11 798.6975 172.25 ;
      END
   END addr1[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 77.82 0.14 77.96 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  915.2425 172.11 915.3825 172.25 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 78.055 0.14 78.195 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  909.045 172.11 909.185 172.25 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  158.4325 172.11 158.5725 172.25 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  159.6075 172.11 159.7475 172.25 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  160.7825 172.11 160.9225 172.25 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  161.9575 172.11 162.0975 172.25 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  163.1325 172.11 163.2725 172.25 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  164.3075 172.11 164.4475 172.25 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  165.4825 172.11 165.6225 172.25 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  166.6575 172.11 166.7975 172.25 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  167.8325 172.11 167.9725 172.25 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  169.0075 172.11 169.1475 172.25 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  170.1825 172.11 170.3225 172.25 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  171.3575 172.11 171.4975 172.25 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  172.5325 172.11 172.6725 172.25 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  173.7075 172.11 173.8475 172.25 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  174.8825 172.11 175.0225 172.25 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  176.0575 172.11 176.1975 172.25 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  177.2325 172.11 177.3725 172.25 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  178.4075 172.11 178.5475 172.25 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  179.5825 172.11 179.7225 172.25 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  180.7575 172.11 180.8975 172.25 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  181.9325 172.11 182.0725 172.25 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  183.1075 172.11 183.2475 172.25 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  184.2825 172.11 184.4225 172.25 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  185.4575 172.11 185.5975 172.25 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  186.6325 172.11 186.7725 172.25 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  187.8075 172.11 187.9475 172.25 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  188.9825 172.11 189.1225 172.25 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  190.1575 172.11 190.2975 172.25 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  191.3325 172.11 191.4725 172.25 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  192.5075 172.11 192.6475 172.25 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  193.6825 172.11 193.8225 172.25 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  194.8575 172.11 194.9975 172.25 ;
      END
   END dout1[31]
   PIN dout1[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  196.0325 172.11 196.1725 172.25 ;
      END
   END dout1[32]
   PIN dout1[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  197.2075 172.11 197.3475 172.25 ;
      END
   END dout1[33]
   PIN dout1[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  198.3825 172.11 198.5225 172.25 ;
      END
   END dout1[34]
   PIN dout1[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  199.5575 172.11 199.6975 172.25 ;
      END
   END dout1[35]
   PIN dout1[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  200.7325 172.11 200.8725 172.25 ;
      END
   END dout1[36]
   PIN dout1[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  201.9075 172.11 202.0475 172.25 ;
      END
   END dout1[37]
   PIN dout1[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  203.0825 172.11 203.2225 172.25 ;
      END
   END dout1[38]
   PIN dout1[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  204.2575 172.11 204.3975 172.25 ;
      END
   END dout1[39]
   PIN dout1[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  205.4325 172.11 205.5725 172.25 ;
      END
   END dout1[40]
   PIN dout1[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  206.6075 172.11 206.7475 172.25 ;
      END
   END dout1[41]
   PIN dout1[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  207.7825 172.11 207.9225 172.25 ;
      END
   END dout1[42]
   PIN dout1[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  208.9575 172.11 209.0975 172.25 ;
      END
   END dout1[43]
   PIN dout1[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  210.1325 172.11 210.2725 172.25 ;
      END
   END dout1[44]
   PIN dout1[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  211.3075 172.11 211.4475 172.25 ;
      END
   END dout1[45]
   PIN dout1[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  212.4825 172.11 212.6225 172.25 ;
      END
   END dout1[46]
   PIN dout1[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  213.6575 172.11 213.7975 172.25 ;
      END
   END dout1[47]
   PIN dout1[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  214.8325 172.11 214.9725 172.25 ;
      END
   END dout1[48]
   PIN dout1[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  216.0075 172.11 216.1475 172.25 ;
      END
   END dout1[49]
   PIN dout1[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  217.1825 172.11 217.3225 172.25 ;
      END
   END dout1[50]
   PIN dout1[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  218.3575 172.11 218.4975 172.25 ;
      END
   END dout1[51]
   PIN dout1[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  219.5325 172.11 219.6725 172.25 ;
      END
   END dout1[52]
   PIN dout1[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  220.7075 172.11 220.8475 172.25 ;
      END
   END dout1[53]
   PIN dout1[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  221.8825 172.11 222.0225 172.25 ;
      END
   END dout1[54]
   PIN dout1[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  223.0575 172.11 223.1975 172.25 ;
      END
   END dout1[55]
   PIN dout1[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  224.2325 172.11 224.3725 172.25 ;
      END
   END dout1[56]
   PIN dout1[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  225.4075 172.11 225.5475 172.25 ;
      END
   END dout1[57]
   PIN dout1[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  226.5825 172.11 226.7225 172.25 ;
      END
   END dout1[58]
   PIN dout1[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  227.7575 172.11 227.8975 172.25 ;
      END
   END dout1[59]
   PIN dout1[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  228.9325 172.11 229.0725 172.25 ;
      END
   END dout1[60]
   PIN dout1[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  230.1075 172.11 230.2475 172.25 ;
      END
   END dout1[61]
   PIN dout1[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  231.2825 172.11 231.4225 172.25 ;
      END
   END dout1[62]
   PIN dout1[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  232.4575 172.11 232.5975 172.25 ;
      END
   END dout1[63]
   PIN dout1[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  233.6325 172.11 233.7725 172.25 ;
      END
   END dout1[64]
   PIN dout1[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  234.8075 172.11 234.9475 172.25 ;
      END
   END dout1[65]
   PIN dout1[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  235.9825 172.11 236.1225 172.25 ;
      END
   END dout1[66]
   PIN dout1[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  237.1575 172.11 237.2975 172.25 ;
      END
   END dout1[67]
   PIN dout1[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  238.3325 172.11 238.4725 172.25 ;
      END
   END dout1[68]
   PIN dout1[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  239.5075 172.11 239.6475 172.25 ;
      END
   END dout1[69]
   PIN dout1[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  240.6825 172.11 240.8225 172.25 ;
      END
   END dout1[70]
   PIN dout1[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  241.8575 172.11 241.9975 172.25 ;
      END
   END dout1[71]
   PIN dout1[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  243.0325 172.11 243.1725 172.25 ;
      END
   END dout1[72]
   PIN dout1[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  244.2075 172.11 244.3475 172.25 ;
      END
   END dout1[73]
   PIN dout1[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  245.3825 172.11 245.5225 172.25 ;
      END
   END dout1[74]
   PIN dout1[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  246.5575 172.11 246.6975 172.25 ;
      END
   END dout1[75]
   PIN dout1[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  247.7325 172.11 247.8725 172.25 ;
      END
   END dout1[76]
   PIN dout1[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  248.9075 172.11 249.0475 172.25 ;
      END
   END dout1[77]
   PIN dout1[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  250.0825 172.11 250.2225 172.25 ;
      END
   END dout1[78]
   PIN dout1[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  251.2575 172.11 251.3975 172.25 ;
      END
   END dout1[79]
   PIN dout1[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  252.4325 172.11 252.5725 172.25 ;
      END
   END dout1[80]
   PIN dout1[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  253.6075 172.11 253.7475 172.25 ;
      END
   END dout1[81]
   PIN dout1[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  254.7825 172.11 254.9225 172.25 ;
      END
   END dout1[82]
   PIN dout1[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  255.9575 172.11 256.0975 172.25 ;
      END
   END dout1[83]
   PIN dout1[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  257.1325 172.11 257.2725 172.25 ;
      END
   END dout1[84]
   PIN dout1[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  258.3075 172.11 258.4475 172.25 ;
      END
   END dout1[85]
   PIN dout1[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  259.4825 172.11 259.6225 172.25 ;
      END
   END dout1[86]
   PIN dout1[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  260.6575 172.11 260.7975 172.25 ;
      END
   END dout1[87]
   PIN dout1[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  261.8325 172.11 261.9725 172.25 ;
      END
   END dout1[88]
   PIN dout1[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  263.0075 172.11 263.1475 172.25 ;
      END
   END dout1[89]
   PIN dout1[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  264.1825 172.11 264.3225 172.25 ;
      END
   END dout1[90]
   PIN dout1[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  265.3575 172.11 265.4975 172.25 ;
      END
   END dout1[91]
   PIN dout1[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  266.5325 172.11 266.6725 172.25 ;
      END
   END dout1[92]
   PIN dout1[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  267.7075 172.11 267.8475 172.25 ;
      END
   END dout1[93]
   PIN dout1[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  268.8825 172.11 269.0225 172.25 ;
      END
   END dout1[94]
   PIN dout1[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  270.0575 172.11 270.1975 172.25 ;
      END
   END dout1[95]
   PIN dout1[96]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  271.2325 172.11 271.3725 172.25 ;
      END
   END dout1[96]
   PIN dout1[97]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  272.4075 172.11 272.5475 172.25 ;
      END
   END dout1[97]
   PIN dout1[98]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  273.5825 172.11 273.7225 172.25 ;
      END
   END dout1[98]
   PIN dout1[99]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  274.7575 172.11 274.8975 172.25 ;
      END
   END dout1[99]
   PIN dout1[100]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  275.9325 172.11 276.0725 172.25 ;
      END
   END dout1[100]
   PIN dout1[101]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  277.1075 172.11 277.2475 172.25 ;
      END
   END dout1[101]
   PIN dout1[102]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  278.2825 172.11 278.4225 172.25 ;
      END
   END dout1[102]
   PIN dout1[103]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  279.4575 172.11 279.5975 172.25 ;
      END
   END dout1[103]
   PIN dout1[104]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  280.6325 172.11 280.7725 172.25 ;
      END
   END dout1[104]
   PIN dout1[105]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  281.8075 172.11 281.9475 172.25 ;
      END
   END dout1[105]
   PIN dout1[106]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  282.9825 172.11 283.1225 172.25 ;
      END
   END dout1[106]
   PIN dout1[107]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  284.1575 172.11 284.2975 172.25 ;
      END
   END dout1[107]
   PIN dout1[108]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  285.3325 172.11 285.4725 172.25 ;
      END
   END dout1[108]
   PIN dout1[109]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  286.5075 172.11 286.6475 172.25 ;
      END
   END dout1[109]
   PIN dout1[110]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  287.6825 172.11 287.8225 172.25 ;
      END
   END dout1[110]
   PIN dout1[111]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  288.8575 172.11 288.9975 172.25 ;
      END
   END dout1[111]
   PIN dout1[112]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  290.0325 172.11 290.1725 172.25 ;
      END
   END dout1[112]
   PIN dout1[113]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  291.2075 172.11 291.3475 172.25 ;
      END
   END dout1[113]
   PIN dout1[114]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  292.3825 172.11 292.5225 172.25 ;
      END
   END dout1[114]
   PIN dout1[115]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  293.5575 172.11 293.6975 172.25 ;
      END
   END dout1[115]
   PIN dout1[116]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  294.7325 172.11 294.8725 172.25 ;
      END
   END dout1[116]
   PIN dout1[117]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  295.9075 172.11 296.0475 172.25 ;
      END
   END dout1[117]
   PIN dout1[118]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  297.0825 172.11 297.2225 172.25 ;
      END
   END dout1[118]
   PIN dout1[119]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  298.2575 172.11 298.3975 172.25 ;
      END
   END dout1[119]
   PIN dout1[120]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  299.4325 172.11 299.5725 172.25 ;
      END
   END dout1[120]
   PIN dout1[121]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  300.6075 172.11 300.7475 172.25 ;
      END
   END dout1[121]
   PIN dout1[122]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  301.7825 172.11 301.9225 172.25 ;
      END
   END dout1[122]
   PIN dout1[123]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  302.9575 172.11 303.0975 172.25 ;
      END
   END dout1[123]
   PIN dout1[124]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  304.1325 172.11 304.2725 172.25 ;
      END
   END dout1[124]
   PIN dout1[125]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  305.3075 172.11 305.4475 172.25 ;
      END
   END dout1[125]
   PIN dout1[126]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  306.4825 172.11 306.6225 172.25 ;
      END
   END dout1[126]
   PIN dout1[127]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  307.6575 172.11 307.7975 172.25 ;
      END
   END dout1[127]
   PIN dout1[128]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  308.8325 172.11 308.9725 172.25 ;
      END
   END dout1[128]
   PIN dout1[129]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  310.0075 172.11 310.1475 172.25 ;
      END
   END dout1[129]
   PIN dout1[130]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  311.1825 172.11 311.3225 172.25 ;
      END
   END dout1[130]
   PIN dout1[131]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  312.3575 172.11 312.4975 172.25 ;
      END
   END dout1[131]
   PIN dout1[132]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  313.5325 172.11 313.6725 172.25 ;
      END
   END dout1[132]
   PIN dout1[133]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  314.7075 172.11 314.8475 172.25 ;
      END
   END dout1[133]
   PIN dout1[134]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  315.8825 172.11 316.0225 172.25 ;
      END
   END dout1[134]
   PIN dout1[135]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  317.0575 172.11 317.1975 172.25 ;
      END
   END dout1[135]
   PIN dout1[136]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  318.2325 172.11 318.3725 172.25 ;
      END
   END dout1[136]
   PIN dout1[137]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  319.4075 172.11 319.5475 172.25 ;
      END
   END dout1[137]
   PIN dout1[138]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  320.5825 172.11 320.7225 172.25 ;
      END
   END dout1[138]
   PIN dout1[139]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  321.7575 172.11 321.8975 172.25 ;
      END
   END dout1[139]
   PIN dout1[140]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  322.9325 172.11 323.0725 172.25 ;
      END
   END dout1[140]
   PIN dout1[141]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  324.1075 172.11 324.2475 172.25 ;
      END
   END dout1[141]
   PIN dout1[142]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  325.2825 172.11 325.4225 172.25 ;
      END
   END dout1[142]
   PIN dout1[143]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  326.4575 172.11 326.5975 172.25 ;
      END
   END dout1[143]
   PIN dout1[144]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  327.6325 172.11 327.7725 172.25 ;
      END
   END dout1[144]
   PIN dout1[145]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  328.8075 172.11 328.9475 172.25 ;
      END
   END dout1[145]
   PIN dout1[146]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  329.9825 172.11 330.1225 172.25 ;
      END
   END dout1[146]
   PIN dout1[147]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  331.1575 172.11 331.2975 172.25 ;
      END
   END dout1[147]
   PIN dout1[148]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  332.3325 172.11 332.4725 172.25 ;
      END
   END dout1[148]
   PIN dout1[149]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  333.5075 172.11 333.6475 172.25 ;
      END
   END dout1[149]
   PIN dout1[150]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  334.6825 172.11 334.8225 172.25 ;
      END
   END dout1[150]
   PIN dout1[151]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  335.8575 172.11 335.9975 172.25 ;
      END
   END dout1[151]
   PIN dout1[152]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  337.0325 172.11 337.1725 172.25 ;
      END
   END dout1[152]
   PIN dout1[153]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  338.2075 172.11 338.3475 172.25 ;
      END
   END dout1[153]
   PIN dout1[154]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  339.3825 172.11 339.5225 172.25 ;
      END
   END dout1[154]
   PIN dout1[155]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  340.5575 172.11 340.6975 172.25 ;
      END
   END dout1[155]
   PIN dout1[156]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  341.7325 172.11 341.8725 172.25 ;
      END
   END dout1[156]
   PIN dout1[157]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  342.9075 172.11 343.0475 172.25 ;
      END
   END dout1[157]
   PIN dout1[158]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  344.0825 172.11 344.2225 172.25 ;
      END
   END dout1[158]
   PIN dout1[159]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  345.2575 172.11 345.3975 172.25 ;
      END
   END dout1[159]
   PIN dout1[160]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  346.4325 172.11 346.5725 172.25 ;
      END
   END dout1[160]
   PIN dout1[161]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  347.6075 172.11 347.7475 172.25 ;
      END
   END dout1[161]
   PIN dout1[162]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  348.7825 172.11 348.9225 172.25 ;
      END
   END dout1[162]
   PIN dout1[163]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  349.9575 172.11 350.0975 172.25 ;
      END
   END dout1[163]
   PIN dout1[164]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  351.1325 172.11 351.2725 172.25 ;
      END
   END dout1[164]
   PIN dout1[165]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  352.3075 172.11 352.4475 172.25 ;
      END
   END dout1[165]
   PIN dout1[166]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  353.4825 172.11 353.6225 172.25 ;
      END
   END dout1[166]
   PIN dout1[167]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  354.6575 172.11 354.7975 172.25 ;
      END
   END dout1[167]
   PIN dout1[168]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  355.8325 172.11 355.9725 172.25 ;
      END
   END dout1[168]
   PIN dout1[169]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  357.0075 172.11 357.1475 172.25 ;
      END
   END dout1[169]
   PIN dout1[170]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  358.1825 172.11 358.3225 172.25 ;
      END
   END dout1[170]
   PIN dout1[171]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  359.3575 172.11 359.4975 172.25 ;
      END
   END dout1[171]
   PIN dout1[172]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  360.5325 172.11 360.6725 172.25 ;
      END
   END dout1[172]
   PIN dout1[173]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  361.7075 172.11 361.8475 172.25 ;
      END
   END dout1[173]
   PIN dout1[174]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  362.8825 172.11 363.0225 172.25 ;
      END
   END dout1[174]
   PIN dout1[175]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  364.0575 172.11 364.1975 172.25 ;
      END
   END dout1[175]
   PIN dout1[176]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  365.2325 172.11 365.3725 172.25 ;
      END
   END dout1[176]
   PIN dout1[177]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  366.4075 172.11 366.5475 172.25 ;
      END
   END dout1[177]
   PIN dout1[178]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  367.5825 172.11 367.7225 172.25 ;
      END
   END dout1[178]
   PIN dout1[179]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  368.7575 172.11 368.8975 172.25 ;
      END
   END dout1[179]
   PIN dout1[180]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  369.9325 172.11 370.0725 172.25 ;
      END
   END dout1[180]
   PIN dout1[181]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  371.1075 172.11 371.2475 172.25 ;
      END
   END dout1[181]
   PIN dout1[182]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  372.2825 172.11 372.4225 172.25 ;
      END
   END dout1[182]
   PIN dout1[183]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  373.4575 172.11 373.5975 172.25 ;
      END
   END dout1[183]
   PIN dout1[184]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  374.6325 172.11 374.7725 172.25 ;
      END
   END dout1[184]
   PIN dout1[185]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  375.8075 172.11 375.9475 172.25 ;
      END
   END dout1[185]
   PIN dout1[186]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  376.9825 172.11 377.1225 172.25 ;
      END
   END dout1[186]
   PIN dout1[187]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  378.1575 172.11 378.2975 172.25 ;
      END
   END dout1[187]
   PIN dout1[188]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  379.3325 172.11 379.4725 172.25 ;
      END
   END dout1[188]
   PIN dout1[189]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  380.5075 172.11 380.6475 172.25 ;
      END
   END dout1[189]
   PIN dout1[190]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  381.6825 172.11 381.8225 172.25 ;
      END
   END dout1[190]
   PIN dout1[191]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  382.8575 172.11 382.9975 172.25 ;
      END
   END dout1[191]
   PIN dout1[192]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  384.0325 172.11 384.1725 172.25 ;
      END
   END dout1[192]
   PIN dout1[193]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  385.2075 172.11 385.3475 172.25 ;
      END
   END dout1[193]
   PIN dout1[194]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  386.3825 172.11 386.5225 172.25 ;
      END
   END dout1[194]
   PIN dout1[195]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  387.5575 172.11 387.6975 172.25 ;
      END
   END dout1[195]
   PIN dout1[196]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  388.7325 172.11 388.8725 172.25 ;
      END
   END dout1[196]
   PIN dout1[197]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  389.9075 172.11 390.0475 172.25 ;
      END
   END dout1[197]
   PIN dout1[198]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  391.0825 172.11 391.2225 172.25 ;
      END
   END dout1[198]
   PIN dout1[199]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  392.2575 172.11 392.3975 172.25 ;
      END
   END dout1[199]
   PIN dout1[200]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  393.4325 172.11 393.5725 172.25 ;
      END
   END dout1[200]
   PIN dout1[201]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  394.6075 172.11 394.7475 172.25 ;
      END
   END dout1[201]
   PIN dout1[202]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  395.7825 172.11 395.9225 172.25 ;
      END
   END dout1[202]
   PIN dout1[203]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  396.9575 172.11 397.0975 172.25 ;
      END
   END dout1[203]
   PIN dout1[204]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  398.1325 172.11 398.2725 172.25 ;
      END
   END dout1[204]
   PIN dout1[205]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  399.3075 172.11 399.4475 172.25 ;
      END
   END dout1[205]
   PIN dout1[206]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  400.4825 172.11 400.6225 172.25 ;
      END
   END dout1[206]
   PIN dout1[207]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  401.6575 172.11 401.7975 172.25 ;
      END
   END dout1[207]
   PIN dout1[208]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  402.8325 172.11 402.9725 172.25 ;
      END
   END dout1[208]
   PIN dout1[209]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  404.0075 172.11 404.1475 172.25 ;
      END
   END dout1[209]
   PIN dout1[210]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  405.1825 172.11 405.3225 172.25 ;
      END
   END dout1[210]
   PIN dout1[211]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  406.3575 172.11 406.4975 172.25 ;
      END
   END dout1[211]
   PIN dout1[212]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  407.5325 172.11 407.6725 172.25 ;
      END
   END dout1[212]
   PIN dout1[213]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  408.7075 172.11 408.8475 172.25 ;
      END
   END dout1[213]
   PIN dout1[214]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  409.8825 172.11 410.0225 172.25 ;
      END
   END dout1[214]
   PIN dout1[215]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  411.0575 172.11 411.1975 172.25 ;
      END
   END dout1[215]
   PIN dout1[216]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  412.2325 172.11 412.3725 172.25 ;
      END
   END dout1[216]
   PIN dout1[217]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  413.4075 172.11 413.5475 172.25 ;
      END
   END dout1[217]
   PIN dout1[218]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  414.5825 172.11 414.7225 172.25 ;
      END
   END dout1[218]
   PIN dout1[219]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  415.7575 172.11 415.8975 172.25 ;
      END
   END dout1[219]
   PIN dout1[220]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  416.9325 172.11 417.0725 172.25 ;
      END
   END dout1[220]
   PIN dout1[221]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  418.1075 172.11 418.2475 172.25 ;
      END
   END dout1[221]
   PIN dout1[222]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  419.2825 172.11 419.4225 172.25 ;
      END
   END dout1[222]
   PIN dout1[223]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  420.4575 172.11 420.5975 172.25 ;
      END
   END dout1[223]
   PIN dout1[224]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  421.6325 172.11 421.7725 172.25 ;
      END
   END dout1[224]
   PIN dout1[225]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  422.8075 172.11 422.9475 172.25 ;
      END
   END dout1[225]
   PIN dout1[226]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  423.9825 172.11 424.1225 172.25 ;
      END
   END dout1[226]
   PIN dout1[227]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  425.1575 172.11 425.2975 172.25 ;
      END
   END dout1[227]
   PIN dout1[228]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  426.3325 172.11 426.4725 172.25 ;
      END
   END dout1[228]
   PIN dout1[229]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  427.5075 172.11 427.6475 172.25 ;
      END
   END dout1[229]
   PIN dout1[230]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  428.6825 172.11 428.8225 172.25 ;
      END
   END dout1[230]
   PIN dout1[231]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  429.8575 172.11 429.9975 172.25 ;
      END
   END dout1[231]
   PIN dout1[232]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  431.0325 172.11 431.1725 172.25 ;
      END
   END dout1[232]
   PIN dout1[233]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  432.2075 172.11 432.3475 172.25 ;
      END
   END dout1[233]
   PIN dout1[234]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  433.3825 172.11 433.5225 172.25 ;
      END
   END dout1[234]
   PIN dout1[235]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  434.5575 172.11 434.6975 172.25 ;
      END
   END dout1[235]
   PIN dout1[236]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  435.7325 172.11 435.8725 172.25 ;
      END
   END dout1[236]
   PIN dout1[237]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  436.9075 172.11 437.0475 172.25 ;
      END
   END dout1[237]
   PIN dout1[238]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  438.0825 172.11 438.2225 172.25 ;
      END
   END dout1[238]
   PIN dout1[239]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  439.2575 172.11 439.3975 172.25 ;
      END
   END dout1[239]
   PIN dout1[240]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  440.4325 172.11 440.5725 172.25 ;
      END
   END dout1[240]
   PIN dout1[241]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  441.6075 172.11 441.7475 172.25 ;
      END
   END dout1[241]
   PIN dout1[242]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  442.7825 172.11 442.9225 172.25 ;
      END
   END dout1[242]
   PIN dout1[243]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  443.9575 172.11 444.0975 172.25 ;
      END
   END dout1[243]
   PIN dout1[244]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  445.1325 172.11 445.2725 172.25 ;
      END
   END dout1[244]
   PIN dout1[245]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  446.3075 172.11 446.4475 172.25 ;
      END
   END dout1[245]
   PIN dout1[246]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  447.4825 172.11 447.6225 172.25 ;
      END
   END dout1[246]
   PIN dout1[247]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  448.6575 172.11 448.7975 172.25 ;
      END
   END dout1[247]
   PIN dout1[248]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  449.8325 172.11 449.9725 172.25 ;
      END
   END dout1[248]
   PIN dout1[249]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  451.0075 172.11 451.1475 172.25 ;
      END
   END dout1[249]
   PIN dout1[250]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  452.1825 172.11 452.3225 172.25 ;
      END
   END dout1[250]
   PIN dout1[251]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  453.3575 172.11 453.4975 172.25 ;
      END
   END dout1[251]
   PIN dout1[252]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  454.5325 172.11 454.6725 172.25 ;
      END
   END dout1[252]
   PIN dout1[253]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  455.7075 172.11 455.8475 172.25 ;
      END
   END dout1[253]
   PIN dout1[254]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  456.8825 172.11 457.0225 172.25 ;
      END
   END dout1[254]
   PIN dout1[255]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  458.0575 172.11 458.1975 172.25 ;
      END
   END dout1[255]
   PIN dout1[256]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  459.2325 172.11 459.3725 172.25 ;
      END
   END dout1[256]
   PIN dout1[257]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  460.4075 172.11 460.5475 172.25 ;
      END
   END dout1[257]
   PIN dout1[258]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  461.5825 172.11 461.7225 172.25 ;
      END
   END dout1[258]
   PIN dout1[259]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  462.7575 172.11 462.8975 172.25 ;
      END
   END dout1[259]
   PIN dout1[260]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  463.9325 172.11 464.0725 172.25 ;
      END
   END dout1[260]
   PIN dout1[261]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  465.1075 172.11 465.2475 172.25 ;
      END
   END dout1[261]
   PIN dout1[262]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  466.2825 172.11 466.4225 172.25 ;
      END
   END dout1[262]
   PIN dout1[263]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  467.4575 172.11 467.5975 172.25 ;
      END
   END dout1[263]
   PIN dout1[264]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  468.6325 172.11 468.7725 172.25 ;
      END
   END dout1[264]
   PIN dout1[265]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  469.8075 172.11 469.9475 172.25 ;
      END
   END dout1[265]
   PIN dout1[266]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  470.9825 172.11 471.1225 172.25 ;
      END
   END dout1[266]
   PIN dout1[267]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  472.1575 172.11 472.2975 172.25 ;
      END
   END dout1[267]
   PIN dout1[268]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  473.3325 172.11 473.4725 172.25 ;
      END
   END dout1[268]
   PIN dout1[269]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  474.5075 172.11 474.6475 172.25 ;
      END
   END dout1[269]
   PIN dout1[270]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  475.6825 172.11 475.8225 172.25 ;
      END
   END dout1[270]
   PIN dout1[271]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  476.8575 172.11 476.9975 172.25 ;
      END
   END dout1[271]
   PIN dout1[272]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  478.0325 172.11 478.1725 172.25 ;
      END
   END dout1[272]
   PIN dout1[273]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  479.2075 172.11 479.3475 172.25 ;
      END
   END dout1[273]
   PIN dout1[274]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  480.3825 172.11 480.5225 172.25 ;
      END
   END dout1[274]
   PIN dout1[275]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  481.5575 172.11 481.6975 172.25 ;
      END
   END dout1[275]
   PIN dout1[276]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  482.7325 172.11 482.8725 172.25 ;
      END
   END dout1[276]
   PIN dout1[277]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  483.9075 172.11 484.0475 172.25 ;
      END
   END dout1[277]
   PIN dout1[278]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  485.0825 172.11 485.2225 172.25 ;
      END
   END dout1[278]
   PIN dout1[279]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  486.2575 172.11 486.3975 172.25 ;
      END
   END dout1[279]
   PIN dout1[280]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  487.4325 172.11 487.5725 172.25 ;
      END
   END dout1[280]
   PIN dout1[281]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  488.6075 172.11 488.7475 172.25 ;
      END
   END dout1[281]
   PIN dout1[282]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  489.7825 172.11 489.9225 172.25 ;
      END
   END dout1[282]
   PIN dout1[283]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  490.9575 172.11 491.0975 172.25 ;
      END
   END dout1[283]
   PIN dout1[284]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  492.1325 172.11 492.2725 172.25 ;
      END
   END dout1[284]
   PIN dout1[285]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  493.3075 172.11 493.4475 172.25 ;
      END
   END dout1[285]
   PIN dout1[286]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  494.4825 172.11 494.6225 172.25 ;
      END
   END dout1[286]
   PIN dout1[287]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  495.6575 172.11 495.7975 172.25 ;
      END
   END dout1[287]
   PIN dout1[288]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  496.8325 172.11 496.9725 172.25 ;
      END
   END dout1[288]
   PIN dout1[289]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  498.0075 172.11 498.1475 172.25 ;
      END
   END dout1[289]
   PIN dout1[290]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  499.1825 172.11 499.3225 172.25 ;
      END
   END dout1[290]
   PIN dout1[291]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  500.3575 172.11 500.4975 172.25 ;
      END
   END dout1[291]
   PIN dout1[292]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  501.5325 172.11 501.6725 172.25 ;
      END
   END dout1[292]
   PIN dout1[293]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  502.7075 172.11 502.8475 172.25 ;
      END
   END dout1[293]
   PIN dout1[294]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  503.8825 172.11 504.0225 172.25 ;
      END
   END dout1[294]
   PIN dout1[295]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  505.0575 172.11 505.1975 172.25 ;
      END
   END dout1[295]
   PIN dout1[296]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  506.2325 172.11 506.3725 172.25 ;
      END
   END dout1[296]
   PIN dout1[297]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  507.4075 172.11 507.5475 172.25 ;
      END
   END dout1[297]
   PIN dout1[298]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  508.5825 172.11 508.7225 172.25 ;
      END
   END dout1[298]
   PIN dout1[299]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  509.7575 172.11 509.8975 172.25 ;
      END
   END dout1[299]
   PIN dout1[300]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  510.9325 172.11 511.0725 172.25 ;
      END
   END dout1[300]
   PIN dout1[301]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  512.1075 172.11 512.2475 172.25 ;
      END
   END dout1[301]
   PIN dout1[302]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  513.2825 172.11 513.4225 172.25 ;
      END
   END dout1[302]
   PIN dout1[303]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  514.4575 172.11 514.5975 172.25 ;
      END
   END dout1[303]
   PIN dout1[304]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  515.6325 172.11 515.7725 172.25 ;
      END
   END dout1[304]
   PIN dout1[305]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  516.8075 172.11 516.9475 172.25 ;
      END
   END dout1[305]
   PIN dout1[306]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  517.9825 172.11 518.1225 172.25 ;
      END
   END dout1[306]
   PIN dout1[307]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  519.1575 172.11 519.2975 172.25 ;
      END
   END dout1[307]
   PIN dout1[308]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  520.3325 172.11 520.4725 172.25 ;
      END
   END dout1[308]
   PIN dout1[309]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  521.5075 172.11 521.6475 172.25 ;
      END
   END dout1[309]
   PIN dout1[310]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  522.6825 172.11 522.8225 172.25 ;
      END
   END dout1[310]
   PIN dout1[311]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  523.8575 172.11 523.9975 172.25 ;
      END
   END dout1[311]
   PIN dout1[312]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  525.0325 172.11 525.1725 172.25 ;
      END
   END dout1[312]
   PIN dout1[313]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  526.2075 172.11 526.3475 172.25 ;
      END
   END dout1[313]
   PIN dout1[314]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  527.3825 172.11 527.5225 172.25 ;
      END
   END dout1[314]
   PIN dout1[315]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  528.5575 172.11 528.6975 172.25 ;
      END
   END dout1[315]
   PIN dout1[316]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  529.7325 172.11 529.8725 172.25 ;
      END
   END dout1[316]
   PIN dout1[317]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  530.9075 172.11 531.0475 172.25 ;
      END
   END dout1[317]
   PIN dout1[318]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  532.0825 172.11 532.2225 172.25 ;
      END
   END dout1[318]
   PIN dout1[319]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  533.2575 172.11 533.3975 172.25 ;
      END
   END dout1[319]
   PIN dout1[320]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  534.4325 172.11 534.5725 172.25 ;
      END
   END dout1[320]
   PIN dout1[321]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  535.6075 172.11 535.7475 172.25 ;
      END
   END dout1[321]
   PIN dout1[322]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  536.7825 172.11 536.9225 172.25 ;
      END
   END dout1[322]
   PIN dout1[323]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  537.9575 172.11 538.0975 172.25 ;
      END
   END dout1[323]
   PIN dout1[324]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  539.1325 172.11 539.2725 172.25 ;
      END
   END dout1[324]
   PIN dout1[325]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  540.3075 172.11 540.4475 172.25 ;
      END
   END dout1[325]
   PIN dout1[326]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  541.4825 172.11 541.6225 172.25 ;
      END
   END dout1[326]
   PIN dout1[327]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  542.6575 172.11 542.7975 172.25 ;
      END
   END dout1[327]
   PIN dout1[328]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  543.8325 172.11 543.9725 172.25 ;
      END
   END dout1[328]
   PIN dout1[329]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  545.0075 172.11 545.1475 172.25 ;
      END
   END dout1[329]
   PIN dout1[330]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  546.1825 172.11 546.3225 172.25 ;
      END
   END dout1[330]
   PIN dout1[331]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  547.3575 172.11 547.4975 172.25 ;
      END
   END dout1[331]
   PIN dout1[332]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  548.5325 172.11 548.6725 172.25 ;
      END
   END dout1[332]
   PIN dout1[333]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  549.7075 172.11 549.8475 172.25 ;
      END
   END dout1[333]
   PIN dout1[334]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  550.8825 172.11 551.0225 172.25 ;
      END
   END dout1[334]
   PIN dout1[335]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  552.0575 172.11 552.1975 172.25 ;
      END
   END dout1[335]
   PIN dout1[336]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  553.2325 172.11 553.3725 172.25 ;
      END
   END dout1[336]
   PIN dout1[337]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  554.4075 172.11 554.5475 172.25 ;
      END
   END dout1[337]
   PIN dout1[338]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  555.5825 172.11 555.7225 172.25 ;
      END
   END dout1[338]
   PIN dout1[339]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  556.7575 172.11 556.8975 172.25 ;
      END
   END dout1[339]
   PIN dout1[340]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  557.9325 172.11 558.0725 172.25 ;
      END
   END dout1[340]
   PIN dout1[341]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  559.1075 172.11 559.2475 172.25 ;
      END
   END dout1[341]
   PIN dout1[342]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  560.2825 172.11 560.4225 172.25 ;
      END
   END dout1[342]
   PIN dout1[343]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  561.4575 172.11 561.5975 172.25 ;
      END
   END dout1[343]
   PIN dout1[344]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  562.6325 172.11 562.7725 172.25 ;
      END
   END dout1[344]
   PIN dout1[345]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  563.8075 172.11 563.9475 172.25 ;
      END
   END dout1[345]
   PIN dout1[346]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  564.9825 172.11 565.1225 172.25 ;
      END
   END dout1[346]
   PIN dout1[347]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  566.1575 172.11 566.2975 172.25 ;
      END
   END dout1[347]
   PIN dout1[348]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  567.3325 172.11 567.4725 172.25 ;
      END
   END dout1[348]
   PIN dout1[349]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  568.5075 172.11 568.6475 172.25 ;
      END
   END dout1[349]
   PIN dout1[350]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  569.6825 172.11 569.8225 172.25 ;
      END
   END dout1[350]
   PIN dout1[351]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  570.8575 172.11 570.9975 172.25 ;
      END
   END dout1[351]
   PIN dout1[352]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  572.0325 172.11 572.1725 172.25 ;
      END
   END dout1[352]
   PIN dout1[353]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  573.2075 172.11 573.3475 172.25 ;
      END
   END dout1[353]
   PIN dout1[354]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  574.3825 172.11 574.5225 172.25 ;
      END
   END dout1[354]
   PIN dout1[355]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  575.5575 172.11 575.6975 172.25 ;
      END
   END dout1[355]
   PIN dout1[356]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  576.7325 172.11 576.8725 172.25 ;
      END
   END dout1[356]
   PIN dout1[357]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  577.9075 172.11 578.0475 172.25 ;
      END
   END dout1[357]
   PIN dout1[358]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  579.0825 172.11 579.2225 172.25 ;
      END
   END dout1[358]
   PIN dout1[359]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  580.2575 172.11 580.3975 172.25 ;
      END
   END dout1[359]
   PIN dout1[360]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  581.4325 172.11 581.5725 172.25 ;
      END
   END dout1[360]
   PIN dout1[361]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  582.6075 172.11 582.7475 172.25 ;
      END
   END dout1[361]
   PIN dout1[362]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  583.7825 172.11 583.9225 172.25 ;
      END
   END dout1[362]
   PIN dout1[363]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  584.9575 172.11 585.0975 172.25 ;
      END
   END dout1[363]
   PIN dout1[364]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  586.1325 172.11 586.2725 172.25 ;
      END
   END dout1[364]
   PIN dout1[365]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  587.3075 172.11 587.4475 172.25 ;
      END
   END dout1[365]
   PIN dout1[366]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  588.4825 172.11 588.6225 172.25 ;
      END
   END dout1[366]
   PIN dout1[367]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  589.6575 172.11 589.7975 172.25 ;
      END
   END dout1[367]
   PIN dout1[368]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  590.8325 172.11 590.9725 172.25 ;
      END
   END dout1[368]
   PIN dout1[369]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  592.0075 172.11 592.1475 172.25 ;
      END
   END dout1[369]
   PIN dout1[370]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  593.1825 172.11 593.3225 172.25 ;
      END
   END dout1[370]
   PIN dout1[371]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  594.3575 172.11 594.4975 172.25 ;
      END
   END dout1[371]
   PIN dout1[372]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  595.5325 172.11 595.6725 172.25 ;
      END
   END dout1[372]
   PIN dout1[373]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  596.7075 172.11 596.8475 172.25 ;
      END
   END dout1[373]
   PIN dout1[374]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  597.8825 172.11 598.0225 172.25 ;
      END
   END dout1[374]
   PIN dout1[375]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  599.0575 172.11 599.1975 172.25 ;
      END
   END dout1[375]
   PIN dout1[376]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  600.2325 172.11 600.3725 172.25 ;
      END
   END dout1[376]
   PIN dout1[377]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  601.4075 172.11 601.5475 172.25 ;
      END
   END dout1[377]
   PIN dout1[378]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  602.5825 172.11 602.7225 172.25 ;
      END
   END dout1[378]
   PIN dout1[379]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  603.7575 172.11 603.8975 172.25 ;
      END
   END dout1[379]
   PIN dout1[380]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  604.9325 172.11 605.0725 172.25 ;
      END
   END dout1[380]
   PIN dout1[381]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  606.1075 172.11 606.2475 172.25 ;
      END
   END dout1[381]
   PIN dout1[382]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  607.2825 172.11 607.4225 172.25 ;
      END
   END dout1[382]
   PIN dout1[383]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  608.4575 172.11 608.5975 172.25 ;
      END
   END dout1[383]
   PIN dout1[384]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  609.6325 172.11 609.7725 172.25 ;
      END
   END dout1[384]
   PIN dout1[385]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  610.8075 172.11 610.9475 172.25 ;
      END
   END dout1[385]
   PIN dout1[386]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  611.9825 172.11 612.1225 172.25 ;
      END
   END dout1[386]
   PIN dout1[387]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  613.1575 172.11 613.2975 172.25 ;
      END
   END dout1[387]
   PIN dout1[388]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  614.3325 172.11 614.4725 172.25 ;
      END
   END dout1[388]
   PIN dout1[389]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  615.5075 172.11 615.6475 172.25 ;
      END
   END dout1[389]
   PIN dout1[390]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  616.6825 172.11 616.8225 172.25 ;
      END
   END dout1[390]
   PIN dout1[391]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  617.8575 172.11 617.9975 172.25 ;
      END
   END dout1[391]
   PIN dout1[392]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  619.0325 172.11 619.1725 172.25 ;
      END
   END dout1[392]
   PIN dout1[393]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  620.2075 172.11 620.3475 172.25 ;
      END
   END dout1[393]
   PIN dout1[394]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  621.3825 172.11 621.5225 172.25 ;
      END
   END dout1[394]
   PIN dout1[395]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  622.5575 172.11 622.6975 172.25 ;
      END
   END dout1[395]
   PIN dout1[396]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  623.7325 172.11 623.8725 172.25 ;
      END
   END dout1[396]
   PIN dout1[397]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  624.9075 172.11 625.0475 172.25 ;
      END
   END dout1[397]
   PIN dout1[398]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  626.0825 172.11 626.2225 172.25 ;
      END
   END dout1[398]
   PIN dout1[399]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  627.2575 172.11 627.3975 172.25 ;
      END
   END dout1[399]
   PIN dout1[400]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  628.4325 172.11 628.5725 172.25 ;
      END
   END dout1[400]
   PIN dout1[401]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  629.6075 172.11 629.7475 172.25 ;
      END
   END dout1[401]
   PIN dout1[402]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  630.7825 172.11 630.9225 172.25 ;
      END
   END dout1[402]
   PIN dout1[403]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  631.9575 172.11 632.0975 172.25 ;
      END
   END dout1[403]
   PIN dout1[404]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  633.1325 172.11 633.2725 172.25 ;
      END
   END dout1[404]
   PIN dout1[405]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  634.3075 172.11 634.4475 172.25 ;
      END
   END dout1[405]
   PIN dout1[406]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  635.4825 172.11 635.6225 172.25 ;
      END
   END dout1[406]
   PIN dout1[407]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  636.6575 172.11 636.7975 172.25 ;
      END
   END dout1[407]
   PIN dout1[408]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  637.8325 172.11 637.9725 172.25 ;
      END
   END dout1[408]
   PIN dout1[409]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  639.0075 172.11 639.1475 172.25 ;
      END
   END dout1[409]
   PIN dout1[410]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  640.1825 172.11 640.3225 172.25 ;
      END
   END dout1[410]
   PIN dout1[411]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  641.3575 172.11 641.4975 172.25 ;
      END
   END dout1[411]
   PIN dout1[412]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  642.5325 172.11 642.6725 172.25 ;
      END
   END dout1[412]
   PIN dout1[413]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  643.7075 172.11 643.8475 172.25 ;
      END
   END dout1[413]
   PIN dout1[414]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  644.8825 172.11 645.0225 172.25 ;
      END
   END dout1[414]
   PIN dout1[415]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  646.0575 172.11 646.1975 172.25 ;
      END
   END dout1[415]
   PIN dout1[416]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  647.2325 172.11 647.3725 172.25 ;
      END
   END dout1[416]
   PIN dout1[417]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  648.4075 172.11 648.5475 172.25 ;
      END
   END dout1[417]
   PIN dout1[418]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  649.5825 172.11 649.7225 172.25 ;
      END
   END dout1[418]
   PIN dout1[419]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  650.7575 172.11 650.8975 172.25 ;
      END
   END dout1[419]
   PIN dout1[420]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  651.9325 172.11 652.0725 172.25 ;
      END
   END dout1[420]
   PIN dout1[421]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  653.1075 172.11 653.2475 172.25 ;
      END
   END dout1[421]
   PIN dout1[422]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  654.2825 172.11 654.4225 172.25 ;
      END
   END dout1[422]
   PIN dout1[423]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  655.4575 172.11 655.5975 172.25 ;
      END
   END dout1[423]
   PIN dout1[424]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  656.6325 172.11 656.7725 172.25 ;
      END
   END dout1[424]
   PIN dout1[425]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  657.8075 172.11 657.9475 172.25 ;
      END
   END dout1[425]
   PIN dout1[426]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  658.9825 172.11 659.1225 172.25 ;
      END
   END dout1[426]
   PIN dout1[427]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  660.1575 172.11 660.2975 172.25 ;
      END
   END dout1[427]
   PIN dout1[428]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  661.3325 172.11 661.4725 172.25 ;
      END
   END dout1[428]
   PIN dout1[429]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  662.5075 172.11 662.6475 172.25 ;
      END
   END dout1[429]
   PIN dout1[430]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  663.6825 172.11 663.8225 172.25 ;
      END
   END dout1[430]
   PIN dout1[431]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  664.8575 172.11 664.9975 172.25 ;
      END
   END dout1[431]
   PIN dout1[432]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  666.0325 172.11 666.1725 172.25 ;
      END
   END dout1[432]
   PIN dout1[433]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  667.2075 172.11 667.3475 172.25 ;
      END
   END dout1[433]
   PIN dout1[434]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  668.3825 172.11 668.5225 172.25 ;
      END
   END dout1[434]
   PIN dout1[435]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  669.5575 172.11 669.6975 172.25 ;
      END
   END dout1[435]
   PIN dout1[436]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  670.7325 172.11 670.8725 172.25 ;
      END
   END dout1[436]
   PIN dout1[437]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  671.9075 172.11 672.0475 172.25 ;
      END
   END dout1[437]
   PIN dout1[438]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  673.0825 172.11 673.2225 172.25 ;
      END
   END dout1[438]
   PIN dout1[439]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  674.2575 172.11 674.3975 172.25 ;
      END
   END dout1[439]
   PIN dout1[440]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  675.4325 172.11 675.5725 172.25 ;
      END
   END dout1[440]
   PIN dout1[441]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  676.6075 172.11 676.7475 172.25 ;
      END
   END dout1[441]
   PIN dout1[442]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  677.7825 172.11 677.9225 172.25 ;
      END
   END dout1[442]
   PIN dout1[443]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  678.9575 172.11 679.0975 172.25 ;
      END
   END dout1[443]
   PIN dout1[444]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  680.1325 172.11 680.2725 172.25 ;
      END
   END dout1[444]
   PIN dout1[445]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  681.3075 172.11 681.4475 172.25 ;
      END
   END dout1[445]
   PIN dout1[446]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  682.4825 172.11 682.6225 172.25 ;
      END
   END dout1[446]
   PIN dout1[447]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  683.6575 172.11 683.7975 172.25 ;
      END
   END dout1[447]
   PIN dout1[448]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  684.8325 172.11 684.9725 172.25 ;
      END
   END dout1[448]
   PIN dout1[449]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  686.0075 172.11 686.1475 172.25 ;
      END
   END dout1[449]
   PIN dout1[450]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  687.1825 172.11 687.3225 172.25 ;
      END
   END dout1[450]
   PIN dout1[451]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  688.3575 172.11 688.4975 172.25 ;
      END
   END dout1[451]
   PIN dout1[452]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  689.5325 172.11 689.6725 172.25 ;
      END
   END dout1[452]
   PIN dout1[453]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  690.7075 172.11 690.8475 172.25 ;
      END
   END dout1[453]
   PIN dout1[454]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  691.8825 172.11 692.0225 172.25 ;
      END
   END dout1[454]
   PIN dout1[455]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  693.0575 172.11 693.1975 172.25 ;
      END
   END dout1[455]
   PIN dout1[456]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  694.2325 172.11 694.3725 172.25 ;
      END
   END dout1[456]
   PIN dout1[457]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  695.4075 172.11 695.5475 172.25 ;
      END
   END dout1[457]
   PIN dout1[458]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  696.5825 172.11 696.7225 172.25 ;
      END
   END dout1[458]
   PIN dout1[459]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  697.7575 172.11 697.8975 172.25 ;
      END
   END dout1[459]
   PIN dout1[460]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  698.9325 172.11 699.0725 172.25 ;
      END
   END dout1[460]
   PIN dout1[461]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  700.1075 172.11 700.2475 172.25 ;
      END
   END dout1[461]
   PIN dout1[462]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  701.2825 172.11 701.4225 172.25 ;
      END
   END dout1[462]
   PIN dout1[463]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  702.4575 172.11 702.5975 172.25 ;
      END
   END dout1[463]
   PIN dout1[464]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  703.6325 172.11 703.7725 172.25 ;
      END
   END dout1[464]
   PIN dout1[465]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  704.8075 172.11 704.9475 172.25 ;
      END
   END dout1[465]
   PIN dout1[466]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  705.9825 172.11 706.1225 172.25 ;
      END
   END dout1[466]
   PIN dout1[467]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  707.1575 172.11 707.2975 172.25 ;
      END
   END dout1[467]
   PIN dout1[468]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  708.3325 172.11 708.4725 172.25 ;
      END
   END dout1[468]
   PIN dout1[469]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  709.5075 172.11 709.6475 172.25 ;
      END
   END dout1[469]
   PIN dout1[470]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  710.6825 172.11 710.8225 172.25 ;
      END
   END dout1[470]
   PIN dout1[471]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  711.8575 172.11 711.9975 172.25 ;
      END
   END dout1[471]
   PIN dout1[472]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  713.0325 172.11 713.1725 172.25 ;
      END
   END dout1[472]
   PIN dout1[473]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  714.2075 172.11 714.3475 172.25 ;
      END
   END dout1[473]
   PIN dout1[474]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  715.3825 172.11 715.5225 172.25 ;
      END
   END dout1[474]
   PIN dout1[475]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  716.5575 172.11 716.6975 172.25 ;
      END
   END dout1[475]
   PIN dout1[476]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  717.7325 172.11 717.8725 172.25 ;
      END
   END dout1[476]
   PIN dout1[477]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  718.9075 172.11 719.0475 172.25 ;
      END
   END dout1[477]
   PIN dout1[478]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  720.0825 172.11 720.2225 172.25 ;
      END
   END dout1[478]
   PIN dout1[479]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  721.2575 172.11 721.3975 172.25 ;
      END
   END dout1[479]
   PIN dout1[480]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  722.4325 172.11 722.5725 172.25 ;
      END
   END dout1[480]
   PIN dout1[481]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  723.6075 172.11 723.7475 172.25 ;
      END
   END dout1[481]
   PIN dout1[482]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  724.7825 172.11 724.9225 172.25 ;
      END
   END dout1[482]
   PIN dout1[483]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  725.9575 172.11 726.0975 172.25 ;
      END
   END dout1[483]
   PIN dout1[484]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  727.1325 172.11 727.2725 172.25 ;
      END
   END dout1[484]
   PIN dout1[485]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  728.3075 172.11 728.4475 172.25 ;
      END
   END dout1[485]
   PIN dout1[486]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  729.4825 172.11 729.6225 172.25 ;
      END
   END dout1[486]
   PIN dout1[487]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  730.6575 172.11 730.7975 172.25 ;
      END
   END dout1[487]
   PIN dout1[488]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  731.8325 172.11 731.9725 172.25 ;
      END
   END dout1[488]
   PIN dout1[489]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  733.0075 172.11 733.1475 172.25 ;
      END
   END dout1[489]
   PIN dout1[490]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  734.1825 172.11 734.3225 172.25 ;
      END
   END dout1[490]
   PIN dout1[491]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  735.3575 172.11 735.4975 172.25 ;
      END
   END dout1[491]
   PIN dout1[492]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  736.5325 172.11 736.6725 172.25 ;
      END
   END dout1[492]
   PIN dout1[493]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  737.7075 172.11 737.8475 172.25 ;
      END
   END dout1[493]
   PIN dout1[494]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  738.8825 172.11 739.0225 172.25 ;
      END
   END dout1[494]
   PIN dout1[495]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  740.0575 172.11 740.1975 172.25 ;
      END
   END dout1[495]
   PIN dout1[496]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  741.2325 172.11 741.3725 172.25 ;
      END
   END dout1[496]
   PIN dout1[497]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  742.4075 172.11 742.5475 172.25 ;
      END
   END dout1[497]
   PIN dout1[498]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  743.5825 172.11 743.7225 172.25 ;
      END
   END dout1[498]
   PIN dout1[499]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  744.7575 172.11 744.8975 172.25 ;
      END
   END dout1[499]
   PIN dout1[500]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  745.9325 172.11 746.0725 172.25 ;
      END
   END dout1[500]
   PIN dout1[501]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  747.1075 172.11 747.2475 172.25 ;
      END
   END dout1[501]
   PIN dout1[502]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  748.2825 172.11 748.4225 172.25 ;
      END
   END dout1[502]
   PIN dout1[503]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  749.4575 172.11 749.5975 172.25 ;
      END
   END dout1[503]
   PIN dout1[504]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  750.6325 172.11 750.7725 172.25 ;
      END
   END dout1[504]
   PIN dout1[505]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  751.8075 172.11 751.9475 172.25 ;
      END
   END dout1[505]
   PIN dout1[506]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  752.9825 172.11 753.1225 172.25 ;
      END
   END dout1[506]
   PIN dout1[507]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  754.1575 172.11 754.2975 172.25 ;
      END
   END dout1[507]
   PIN dout1[508]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  755.3325 172.11 755.4725 172.25 ;
      END
   END dout1[508]
   PIN dout1[509]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  756.5075 172.11 756.6475 172.25 ;
      END
   END dout1[509]
   PIN dout1[510]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  757.6825 172.11 757.8225 172.25 ;
      END
   END dout1[510]
   PIN dout1[511]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  758.8575 172.11 758.9975 172.25 ;
      END
   END dout1[511]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 1589.735 172.11 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 1589.735 172.11 ;
   LAYER  metal3 ;
      RECT  0.14 0.14 0.28 77.68 ;
      RECT  0.28 0.14 1589.735 77.68 ;
      RECT  0.28 77.68 1589.735 78.1 ;
      RECT  0.28 78.1 1589.735 172.11 ;
      RECT  0.14 78.335 0.28 172.11 ;
   LAYER  metal4 ;
      RECT  0.14 0.14 125.4875 0.42 ;
      RECT  125.4875 0.42 126.1875 172.11 ;
      RECT  126.1875 0.14 128.3475 0.42 ;
      RECT  129.0475 0.14 131.2075 0.42 ;
      RECT  131.9075 0.14 134.0675 0.42 ;
      RECT  134.7675 0.14 136.9275 0.42 ;
      RECT  137.6275 0.14 139.7875 0.42 ;
      RECT  140.4875 0.14 142.6475 0.42 ;
      RECT  143.3475 0.14 145.5075 0.42 ;
      RECT  146.2075 0.14 148.3675 0.42 ;
      RECT  149.0675 0.14 151.2275 0.42 ;
      RECT  151.9275 0.14 154.0875 0.42 ;
      RECT  154.7875 0.14 156.9475 0.42 ;
      RECT  157.6475 0.14 159.8075 0.42 ;
      RECT  160.5075 0.14 162.6675 0.42 ;
      RECT  163.3675 0.14 165.5275 0.42 ;
      RECT  166.2275 0.14 168.3875 0.42 ;
      RECT  169.0875 0.14 171.2475 0.42 ;
      RECT  171.9475 0.14 174.1075 0.42 ;
      RECT  174.8075 0.14 176.9675 0.42 ;
      RECT  177.6675 0.14 179.8275 0.42 ;
      RECT  180.5275 0.14 182.6875 0.42 ;
      RECT  183.3875 0.14 185.5475 0.42 ;
      RECT  186.2475 0.14 188.4075 0.42 ;
      RECT  189.1075 0.14 191.2675 0.42 ;
      RECT  191.9675 0.14 194.1275 0.42 ;
      RECT  194.8275 0.14 196.9875 0.42 ;
      RECT  197.6875 0.14 199.8475 0.42 ;
      RECT  200.5475 0.14 202.7075 0.42 ;
      RECT  203.4075 0.14 205.5675 0.42 ;
      RECT  206.2675 0.14 208.4275 0.42 ;
      RECT  209.1275 0.14 211.2875 0.42 ;
      RECT  211.9875 0.14 214.1475 0.42 ;
      RECT  214.8475 0.14 217.0075 0.42 ;
      RECT  217.7075 0.14 219.8675 0.42 ;
      RECT  220.5675 0.14 222.7275 0.42 ;
      RECT  223.4275 0.14 225.5875 0.42 ;
      RECT  226.2875 0.14 228.4475 0.42 ;
      RECT  229.1475 0.14 231.3075 0.42 ;
      RECT  232.0075 0.14 234.1675 0.42 ;
      RECT  234.8675 0.14 237.0275 0.42 ;
      RECT  237.7275 0.14 239.8875 0.42 ;
      RECT  240.5875 0.14 242.7475 0.42 ;
      RECT  243.4475 0.14 245.6075 0.42 ;
      RECT  246.3075 0.14 248.4675 0.42 ;
      RECT  249.1675 0.14 251.3275 0.42 ;
      RECT  252.0275 0.14 254.1875 0.42 ;
      RECT  254.8875 0.14 257.0475 0.42 ;
      RECT  257.7475 0.14 259.9075 0.42 ;
      RECT  260.6075 0.14 262.7675 0.42 ;
      RECT  263.4675 0.14 265.6275 0.42 ;
      RECT  266.3275 0.14 268.4875 0.42 ;
      RECT  269.1875 0.14 271.3475 0.42 ;
      RECT  272.0475 0.14 274.2075 0.42 ;
      RECT  274.9075 0.14 277.0675 0.42 ;
      RECT  277.7675 0.14 279.9275 0.42 ;
      RECT  280.6275 0.14 282.7875 0.42 ;
      RECT  283.4875 0.14 285.6475 0.42 ;
      RECT  286.3475 0.14 288.5075 0.42 ;
      RECT  289.2075 0.14 291.3675 0.42 ;
      RECT  292.0675 0.14 294.2275 0.42 ;
      RECT  294.9275 0.14 297.0875 0.42 ;
      RECT  297.7875 0.14 299.9475 0.42 ;
      RECT  300.6475 0.14 302.8075 0.42 ;
      RECT  303.5075 0.14 305.6675 0.42 ;
      RECT  306.3675 0.14 308.5275 0.42 ;
      RECT  309.2275 0.14 311.3875 0.42 ;
      RECT  312.0875 0.14 314.2475 0.42 ;
      RECT  314.9475 0.14 317.1075 0.42 ;
      RECT  317.8075 0.14 319.9675 0.42 ;
      RECT  320.6675 0.14 322.8275 0.42 ;
      RECT  323.5275 0.14 325.6875 0.42 ;
      RECT  326.3875 0.14 328.5475 0.42 ;
      RECT  329.2475 0.14 331.4075 0.42 ;
      RECT  332.1075 0.14 334.2675 0.42 ;
      RECT  334.9675 0.14 337.1275 0.42 ;
      RECT  337.8275 0.14 339.9875 0.42 ;
      RECT  340.6875 0.14 342.8475 0.42 ;
      RECT  343.5475 0.14 345.7075 0.42 ;
      RECT  346.4075 0.14 348.5675 0.42 ;
      RECT  349.2675 0.14 351.4275 0.42 ;
      RECT  352.1275 0.14 354.2875 0.42 ;
      RECT  354.9875 0.14 357.1475 0.42 ;
      RECT  357.8475 0.14 360.0075 0.42 ;
      RECT  360.7075 0.14 362.8675 0.42 ;
      RECT  363.5675 0.14 365.7275 0.42 ;
      RECT  366.4275 0.14 368.5875 0.42 ;
      RECT  369.2875 0.14 371.4475 0.42 ;
      RECT  372.1475 0.14 374.3075 0.42 ;
      RECT  375.0075 0.14 377.1675 0.42 ;
      RECT  377.8675 0.14 380.0275 0.42 ;
      RECT  380.7275 0.14 382.8875 0.42 ;
      RECT  383.5875 0.14 385.7475 0.42 ;
      RECT  386.4475 0.14 388.6075 0.42 ;
      RECT  389.3075 0.14 391.4675 0.42 ;
      RECT  392.1675 0.14 394.3275 0.42 ;
      RECT  395.0275 0.14 397.1875 0.42 ;
      RECT  397.8875 0.14 400.0475 0.42 ;
      RECT  400.7475 0.14 402.9075 0.42 ;
      RECT  403.6075 0.14 405.7675 0.42 ;
      RECT  406.4675 0.14 408.6275 0.42 ;
      RECT  409.3275 0.14 411.4875 0.42 ;
      RECT  412.1875 0.14 414.3475 0.42 ;
      RECT  415.0475 0.14 417.2075 0.42 ;
      RECT  417.9075 0.14 420.0675 0.42 ;
      RECT  420.7675 0.14 422.9275 0.42 ;
      RECT  423.6275 0.14 425.7875 0.42 ;
      RECT  426.4875 0.14 428.6475 0.42 ;
      RECT  429.3475 0.14 431.5075 0.42 ;
      RECT  432.2075 0.14 434.3675 0.42 ;
      RECT  435.0675 0.14 437.2275 0.42 ;
      RECT  437.9275 0.14 440.0875 0.42 ;
      RECT  440.7875 0.14 442.9475 0.42 ;
      RECT  443.6475 0.14 445.8075 0.42 ;
      RECT  446.5075 0.14 448.6675 0.42 ;
      RECT  449.3675 0.14 451.5275 0.42 ;
      RECT  452.2275 0.14 454.3875 0.42 ;
      RECT  455.0875 0.14 457.2475 0.42 ;
      RECT  457.9475 0.14 460.1075 0.42 ;
      RECT  460.8075 0.14 462.9675 0.42 ;
      RECT  463.6675 0.14 465.8275 0.42 ;
      RECT  466.5275 0.14 468.6875 0.42 ;
      RECT  469.3875 0.14 471.5475 0.42 ;
      RECT  472.2475 0.14 474.4075 0.42 ;
      RECT  475.1075 0.14 477.2675 0.42 ;
      RECT  477.9675 0.14 480.1275 0.42 ;
      RECT  480.8275 0.14 482.9875 0.42 ;
      RECT  483.6875 0.14 485.8475 0.42 ;
      RECT  486.5475 0.14 488.7075 0.42 ;
      RECT  489.4075 0.14 491.5675 0.42 ;
      RECT  492.2675 0.14 494.4275 0.42 ;
      RECT  495.1275 0.14 497.2875 0.42 ;
      RECT  497.9875 0.14 500.1475 0.42 ;
      RECT  500.8475 0.14 503.0075 0.42 ;
      RECT  503.7075 0.14 505.8675 0.42 ;
      RECT  506.5675 0.14 508.7275 0.42 ;
      RECT  509.4275 0.14 511.5875 0.42 ;
      RECT  512.2875 0.14 514.4475 0.42 ;
      RECT  515.1475 0.14 517.3075 0.42 ;
      RECT  518.0075 0.14 520.1675 0.42 ;
      RECT  520.8675 0.14 523.0275 0.42 ;
      RECT  523.7275 0.14 525.8875 0.42 ;
      RECT  526.5875 0.14 528.7475 0.42 ;
      RECT  529.4475 0.14 531.6075 0.42 ;
      RECT  532.3075 0.14 534.4675 0.42 ;
      RECT  535.1675 0.14 537.3275 0.42 ;
      RECT  538.0275 0.14 540.1875 0.42 ;
      RECT  540.8875 0.14 543.0475 0.42 ;
      RECT  543.7475 0.14 545.9075 0.42 ;
      RECT  546.6075 0.14 548.7675 0.42 ;
      RECT  549.4675 0.14 551.6275 0.42 ;
      RECT  552.3275 0.14 554.4875 0.42 ;
      RECT  555.1875 0.14 557.3475 0.42 ;
      RECT  558.0475 0.14 560.2075 0.42 ;
      RECT  560.9075 0.14 563.0675 0.42 ;
      RECT  563.7675 0.14 565.9275 0.42 ;
      RECT  566.6275 0.14 568.7875 0.42 ;
      RECT  569.4875 0.14 571.6475 0.42 ;
      RECT  572.3475 0.14 574.5075 0.42 ;
      RECT  575.2075 0.14 577.3675 0.42 ;
      RECT  578.0675 0.14 580.2275 0.42 ;
      RECT  580.9275 0.14 583.0875 0.42 ;
      RECT  583.7875 0.14 585.9475 0.42 ;
      RECT  586.6475 0.14 588.8075 0.42 ;
      RECT  589.5075 0.14 591.6675 0.42 ;
      RECT  592.3675 0.14 594.5275 0.42 ;
      RECT  595.2275 0.14 597.3875 0.42 ;
      RECT  598.0875 0.14 600.2475 0.42 ;
      RECT  600.9475 0.14 603.1075 0.42 ;
      RECT  603.8075 0.14 605.9675 0.42 ;
      RECT  606.6675 0.14 608.8275 0.42 ;
      RECT  609.5275 0.14 611.6875 0.42 ;
      RECT  612.3875 0.14 614.5475 0.42 ;
      RECT  615.2475 0.14 617.4075 0.42 ;
      RECT  618.1075 0.14 620.2675 0.42 ;
      RECT  620.9675 0.14 623.1275 0.42 ;
      RECT  623.8275 0.14 625.9875 0.42 ;
      RECT  626.6875 0.14 628.8475 0.42 ;
      RECT  629.5475 0.14 631.7075 0.42 ;
      RECT  632.4075 0.14 634.5675 0.42 ;
      RECT  635.2675 0.14 637.4275 0.42 ;
      RECT  638.1275 0.14 640.2875 0.42 ;
      RECT  640.9875 0.14 643.1475 0.42 ;
      RECT  643.8475 0.14 646.0075 0.42 ;
      RECT  646.7075 0.14 648.8675 0.42 ;
      RECT  649.5675 0.14 651.7275 0.42 ;
      RECT  652.4275 0.14 654.5875 0.42 ;
      RECT  655.2875 0.14 657.4475 0.42 ;
      RECT  658.1475 0.14 660.3075 0.42 ;
      RECT  661.0075 0.14 663.1675 0.42 ;
      RECT  663.8675 0.14 666.0275 0.42 ;
      RECT  666.7275 0.14 668.8875 0.42 ;
      RECT  669.5875 0.14 671.7475 0.42 ;
      RECT  672.4475 0.14 674.6075 0.42 ;
      RECT  675.3075 0.14 677.4675 0.42 ;
      RECT  678.1675 0.14 680.3275 0.42 ;
      RECT  681.0275 0.14 683.1875 0.42 ;
      RECT  683.8875 0.14 686.0475 0.42 ;
      RECT  686.7475 0.14 688.9075 0.42 ;
      RECT  689.6075 0.14 691.7675 0.42 ;
      RECT  692.4675 0.14 694.6275 0.42 ;
      RECT  695.3275 0.14 697.4875 0.42 ;
      RECT  698.1875 0.14 700.3475 0.42 ;
      RECT  701.0475 0.14 703.2075 0.42 ;
      RECT  703.9075 0.14 706.0675 0.42 ;
      RECT  706.7675 0.14 708.9275 0.42 ;
      RECT  709.6275 0.14 711.7875 0.42 ;
      RECT  712.4875 0.14 714.6475 0.42 ;
      RECT  715.3475 0.14 717.5075 0.42 ;
      RECT  718.2075 0.14 720.3675 0.42 ;
      RECT  721.0675 0.14 723.2275 0.42 ;
      RECT  723.9275 0.14 726.0875 0.42 ;
      RECT  726.7875 0.14 728.9475 0.42 ;
      RECT  729.6475 0.14 731.8075 0.42 ;
      RECT  732.5075 0.14 734.6675 0.42 ;
      RECT  735.3675 0.14 737.5275 0.42 ;
      RECT  738.2275 0.14 740.3875 0.42 ;
      RECT  741.0875 0.14 743.2475 0.42 ;
      RECT  743.9475 0.14 746.1075 0.42 ;
      RECT  746.8075 0.14 748.9675 0.42 ;
      RECT  749.6675 0.14 751.8275 0.42 ;
      RECT  752.5275 0.14 754.6875 0.42 ;
      RECT  755.3875 0.14 757.5475 0.42 ;
      RECT  758.2475 0.14 760.4075 0.42 ;
      RECT  761.1075 0.14 763.2675 0.42 ;
      RECT  763.9675 0.14 766.1275 0.42 ;
      RECT  766.8275 0.14 768.9875 0.42 ;
      RECT  769.6875 0.14 771.8475 0.42 ;
      RECT  772.5475 0.14 774.7075 0.42 ;
      RECT  775.4075 0.14 777.5675 0.42 ;
      RECT  778.2675 0.14 780.4275 0.42 ;
      RECT  781.1275 0.14 783.2875 0.42 ;
      RECT  783.9875 0.14 786.1475 0.42 ;
      RECT  786.8475 0.14 789.0075 0.42 ;
      RECT  789.7075 0.14 791.8675 0.42 ;
      RECT  792.5675 0.14 794.7275 0.42 ;
      RECT  795.4275 0.14 797.5875 0.42 ;
      RECT  798.2875 0.14 800.4475 0.42 ;
      RECT  801.1475 0.14 803.3075 0.42 ;
      RECT  804.0075 0.14 806.1675 0.42 ;
      RECT  806.8675 0.14 809.0275 0.42 ;
      RECT  809.7275 0.14 811.8875 0.42 ;
      RECT  812.5875 0.14 814.7475 0.42 ;
      RECT  815.4475 0.14 817.6075 0.42 ;
      RECT  818.3075 0.14 820.4675 0.42 ;
      RECT  821.1675 0.14 823.3275 0.42 ;
      RECT  824.0275 0.14 826.1875 0.42 ;
      RECT  826.8875 0.14 829.0475 0.42 ;
      RECT  829.7475 0.14 831.9075 0.42 ;
      RECT  832.6075 0.14 834.7675 0.42 ;
      RECT  835.4675 0.14 837.6275 0.42 ;
      RECT  838.3275 0.14 840.4875 0.42 ;
      RECT  841.1875 0.14 843.3475 0.42 ;
      RECT  844.0475 0.14 846.2075 0.42 ;
      RECT  846.9075 0.14 849.0675 0.42 ;
      RECT  849.7675 0.14 851.9275 0.42 ;
      RECT  852.6275 0.14 854.7875 0.42 ;
      RECT  855.4875 0.14 857.6475 0.42 ;
      RECT  858.3475 0.14 860.5075 0.42 ;
      RECT  861.2075 0.14 863.3675 0.42 ;
      RECT  864.0675 0.14 866.2275 0.42 ;
      RECT  866.9275 0.14 869.0875 0.42 ;
      RECT  869.7875 0.14 871.9475 0.42 ;
      RECT  872.6475 0.14 874.8075 0.42 ;
      RECT  875.5075 0.14 877.6675 0.42 ;
      RECT  878.3675 0.14 880.5275 0.42 ;
      RECT  881.2275 0.14 883.3875 0.42 ;
      RECT  884.0875 0.14 886.2475 0.42 ;
      RECT  886.9475 0.14 889.1075 0.42 ;
      RECT  889.8075 0.14 891.9675 0.42 ;
      RECT  892.6675 0.14 894.8275 0.42 ;
      RECT  895.5275 0.14 897.6875 0.42 ;
      RECT  898.3875 0.14 900.5475 0.42 ;
      RECT  901.2475 0.14 903.4075 0.42 ;
      RECT  904.1075 0.14 906.2675 0.42 ;
      RECT  906.9675 0.14 909.1275 0.42 ;
      RECT  909.8275 0.14 911.9875 0.42 ;
      RECT  912.6875 0.14 914.8475 0.42 ;
      RECT  915.5475 0.14 917.7075 0.42 ;
      RECT  918.4075 0.14 920.5675 0.42 ;
      RECT  921.2675 0.14 923.4275 0.42 ;
      RECT  924.1275 0.14 926.2875 0.42 ;
      RECT  926.9875 0.14 929.1475 0.42 ;
      RECT  929.8475 0.14 932.0075 0.42 ;
      RECT  932.7075 0.14 934.8675 0.42 ;
      RECT  935.5675 0.14 937.7275 0.42 ;
      RECT  938.4275 0.14 940.5875 0.42 ;
      RECT  941.2875 0.14 943.4475 0.42 ;
      RECT  944.1475 0.14 946.3075 0.42 ;
      RECT  947.0075 0.14 949.1675 0.42 ;
      RECT  949.8675 0.14 952.0275 0.42 ;
      RECT  952.7275 0.14 954.8875 0.42 ;
      RECT  955.5875 0.14 957.7475 0.42 ;
      RECT  958.4475 0.14 960.6075 0.42 ;
      RECT  961.3075 0.14 963.4675 0.42 ;
      RECT  964.1675 0.14 966.3275 0.42 ;
      RECT  967.0275 0.14 969.1875 0.42 ;
      RECT  969.8875 0.14 972.0475 0.42 ;
      RECT  972.7475 0.14 974.9075 0.42 ;
      RECT  975.6075 0.14 977.7675 0.42 ;
      RECT  978.4675 0.14 980.6275 0.42 ;
      RECT  981.3275 0.14 983.4875 0.42 ;
      RECT  984.1875 0.14 986.3475 0.42 ;
      RECT  987.0475 0.14 989.2075 0.42 ;
      RECT  989.9075 0.14 992.0675 0.42 ;
      RECT  992.7675 0.14 994.9275 0.42 ;
      RECT  995.6275 0.14 997.7875 0.42 ;
      RECT  998.4875 0.14 1000.6475 0.42 ;
      RECT  1001.3475 0.14 1003.5075 0.42 ;
      RECT  1004.2075 0.14 1006.3675 0.42 ;
      RECT  1007.0675 0.14 1009.2275 0.42 ;
      RECT  1009.9275 0.14 1012.0875 0.42 ;
      RECT  1012.7875 0.14 1014.9475 0.42 ;
      RECT  1015.6475 0.14 1017.8075 0.42 ;
      RECT  1018.5075 0.14 1020.6675 0.42 ;
      RECT  1021.3675 0.14 1023.5275 0.42 ;
      RECT  1024.2275 0.14 1026.3875 0.42 ;
      RECT  1027.0875 0.14 1029.2475 0.42 ;
      RECT  1029.9475 0.14 1032.1075 0.42 ;
      RECT  1032.8075 0.14 1034.9675 0.42 ;
      RECT  1035.6675 0.14 1037.8275 0.42 ;
      RECT  1038.5275 0.14 1040.6875 0.42 ;
      RECT  1041.3875 0.14 1043.5475 0.42 ;
      RECT  1044.2475 0.14 1046.4075 0.42 ;
      RECT  1047.1075 0.14 1049.2675 0.42 ;
      RECT  1049.9675 0.14 1052.1275 0.42 ;
      RECT  1052.8275 0.14 1054.9875 0.42 ;
      RECT  1055.6875 0.14 1057.8475 0.42 ;
      RECT  1058.5475 0.14 1060.7075 0.42 ;
      RECT  1061.4075 0.14 1063.5675 0.42 ;
      RECT  1064.2675 0.14 1066.4275 0.42 ;
      RECT  1067.1275 0.14 1069.2875 0.42 ;
      RECT  1069.9875 0.14 1072.1475 0.42 ;
      RECT  1072.8475 0.14 1075.0075 0.42 ;
      RECT  1075.7075 0.14 1077.8675 0.42 ;
      RECT  1078.5675 0.14 1080.7275 0.42 ;
      RECT  1081.4275 0.14 1083.5875 0.42 ;
      RECT  1084.2875 0.14 1086.4475 0.42 ;
      RECT  1087.1475 0.14 1089.3075 0.42 ;
      RECT  1090.0075 0.14 1092.1675 0.42 ;
      RECT  1092.8675 0.14 1095.0275 0.42 ;
      RECT  1095.7275 0.14 1097.8875 0.42 ;
      RECT  1098.5875 0.14 1100.7475 0.42 ;
      RECT  1101.4475 0.14 1103.6075 0.42 ;
      RECT  1104.3075 0.14 1106.4675 0.42 ;
      RECT  1107.1675 0.14 1109.3275 0.42 ;
      RECT  1110.0275 0.14 1112.1875 0.42 ;
      RECT  1112.8875 0.14 1115.0475 0.42 ;
      RECT  1115.7475 0.14 1117.9075 0.42 ;
      RECT  1118.6075 0.14 1120.7675 0.42 ;
      RECT  1121.4675 0.14 1123.6275 0.42 ;
      RECT  1124.3275 0.14 1126.4875 0.42 ;
      RECT  1127.1875 0.14 1129.3475 0.42 ;
      RECT  1130.0475 0.14 1132.2075 0.42 ;
      RECT  1132.9075 0.14 1135.0675 0.42 ;
      RECT  1135.7675 0.14 1137.9275 0.42 ;
      RECT  1138.6275 0.14 1140.7875 0.42 ;
      RECT  1141.4875 0.14 1143.6475 0.42 ;
      RECT  1144.3475 0.14 1146.5075 0.42 ;
      RECT  1147.2075 0.14 1149.3675 0.42 ;
      RECT  1150.0675 0.14 1152.2275 0.42 ;
      RECT  1152.9275 0.14 1155.0875 0.42 ;
      RECT  1155.7875 0.14 1157.9475 0.42 ;
      RECT  1158.6475 0.14 1160.8075 0.42 ;
      RECT  1161.5075 0.14 1163.6675 0.42 ;
      RECT  1164.3675 0.14 1166.5275 0.42 ;
      RECT  1167.2275 0.14 1169.3875 0.42 ;
      RECT  1170.0875 0.14 1172.2475 0.42 ;
      RECT  1172.9475 0.14 1175.1075 0.42 ;
      RECT  1175.8075 0.14 1177.9675 0.42 ;
      RECT  1178.6675 0.14 1180.8275 0.42 ;
      RECT  1181.5275 0.14 1183.6875 0.42 ;
      RECT  1184.3875 0.14 1186.5475 0.42 ;
      RECT  1187.2475 0.14 1189.4075 0.42 ;
      RECT  1190.1075 0.14 1192.2675 0.42 ;
      RECT  1192.9675 0.14 1195.1275 0.42 ;
      RECT  1195.8275 0.14 1197.9875 0.42 ;
      RECT  1198.6875 0.14 1200.8475 0.42 ;
      RECT  1201.5475 0.14 1203.7075 0.42 ;
      RECT  1204.4075 0.14 1206.5675 0.42 ;
      RECT  1207.2675 0.14 1209.4275 0.42 ;
      RECT  1210.1275 0.14 1212.2875 0.42 ;
      RECT  1212.9875 0.14 1215.1475 0.42 ;
      RECT  1215.8475 0.14 1218.0075 0.42 ;
      RECT  1218.7075 0.14 1220.8675 0.42 ;
      RECT  1221.5675 0.14 1223.7275 0.42 ;
      RECT  1224.4275 0.14 1226.5875 0.42 ;
      RECT  1227.2875 0.14 1229.4475 0.42 ;
      RECT  1230.1475 0.14 1232.3075 0.42 ;
      RECT  1233.0075 0.14 1235.1675 0.42 ;
      RECT  1235.8675 0.14 1238.0275 0.42 ;
      RECT  1238.7275 0.14 1240.8875 0.42 ;
      RECT  1241.5875 0.14 1243.7475 0.42 ;
      RECT  1244.4475 0.14 1246.6075 0.42 ;
      RECT  1247.3075 0.14 1249.4675 0.42 ;
      RECT  1250.1675 0.14 1252.3275 0.42 ;
      RECT  1253.0275 0.14 1255.1875 0.42 ;
      RECT  1255.8875 0.14 1258.0475 0.42 ;
      RECT  1258.7475 0.14 1260.9075 0.42 ;
      RECT  1261.6075 0.14 1263.7675 0.42 ;
      RECT  1264.4675 0.14 1266.6275 0.42 ;
      RECT  1267.3275 0.14 1269.4875 0.42 ;
      RECT  1270.1875 0.14 1272.3475 0.42 ;
      RECT  1273.0475 0.14 1275.2075 0.42 ;
      RECT  1275.9075 0.14 1278.0675 0.42 ;
      RECT  1278.7675 0.14 1280.9275 0.42 ;
      RECT  1281.6275 0.14 1283.7875 0.42 ;
      RECT  1284.4875 0.14 1286.6475 0.42 ;
      RECT  1287.3475 0.14 1289.5075 0.42 ;
      RECT  1290.2075 0.14 1292.3675 0.42 ;
      RECT  1293.0675 0.14 1295.2275 0.42 ;
      RECT  1295.9275 0.14 1298.0875 0.42 ;
      RECT  1298.7875 0.14 1300.9475 0.42 ;
      RECT  1301.6475 0.14 1303.8075 0.42 ;
      RECT  1304.5075 0.14 1306.6675 0.42 ;
      RECT  1307.3675 0.14 1309.5275 0.42 ;
      RECT  1310.2275 0.14 1312.3875 0.42 ;
      RECT  1313.0875 0.14 1315.2475 0.42 ;
      RECT  1315.9475 0.14 1318.1075 0.42 ;
      RECT  1318.8075 0.14 1320.9675 0.42 ;
      RECT  1321.6675 0.14 1323.8275 0.42 ;
      RECT  1324.5275 0.14 1326.6875 0.42 ;
      RECT  1327.3875 0.14 1329.5475 0.42 ;
      RECT  1330.2475 0.14 1332.4075 0.42 ;
      RECT  1333.1075 0.14 1335.2675 0.42 ;
      RECT  1335.9675 0.14 1338.1275 0.42 ;
      RECT  1338.8275 0.14 1340.9875 0.42 ;
      RECT  1341.6875 0.14 1343.8475 0.42 ;
      RECT  1344.5475 0.14 1346.7075 0.42 ;
      RECT  1347.4075 0.14 1349.5675 0.42 ;
      RECT  1350.2675 0.14 1352.4275 0.42 ;
      RECT  1353.1275 0.14 1355.2875 0.42 ;
      RECT  1355.9875 0.14 1358.1475 0.42 ;
      RECT  1358.8475 0.14 1361.0075 0.42 ;
      RECT  1361.7075 0.14 1363.8675 0.42 ;
      RECT  1364.5675 0.14 1366.7275 0.42 ;
      RECT  1367.4275 0.14 1369.5875 0.42 ;
      RECT  1370.2875 0.14 1372.4475 0.42 ;
      RECT  1373.1475 0.14 1375.3075 0.42 ;
      RECT  1376.0075 0.14 1378.1675 0.42 ;
      RECT  1378.8675 0.14 1381.0275 0.42 ;
      RECT  1381.7275 0.14 1383.8875 0.42 ;
      RECT  1384.5875 0.14 1386.7475 0.42 ;
      RECT  1387.4475 0.14 1389.6075 0.42 ;
      RECT  1390.3075 0.14 1392.4675 0.42 ;
      RECT  1393.1675 0.14 1395.3275 0.42 ;
      RECT  1396.0275 0.14 1398.1875 0.42 ;
      RECT  1398.8875 0.14 1401.0475 0.42 ;
      RECT  1401.7475 0.14 1403.9075 0.42 ;
      RECT  1404.6075 0.14 1406.7675 0.42 ;
      RECT  1407.4675 0.14 1409.6275 0.42 ;
      RECT  1410.3275 0.14 1412.4875 0.42 ;
      RECT  1413.1875 0.14 1415.3475 0.42 ;
      RECT  1416.0475 0.14 1418.2075 0.42 ;
      RECT  1418.9075 0.14 1421.0675 0.42 ;
      RECT  1421.7675 0.14 1423.9275 0.42 ;
      RECT  1424.6275 0.14 1426.7875 0.42 ;
      RECT  1427.4875 0.14 1429.6475 0.42 ;
      RECT  1430.3475 0.14 1432.5075 0.42 ;
      RECT  1433.2075 0.14 1435.3675 0.42 ;
      RECT  1436.0675 0.14 1438.2275 0.42 ;
      RECT  1438.9275 0.14 1441.0875 0.42 ;
      RECT  1441.7875 0.14 1443.9475 0.42 ;
      RECT  1444.6475 0.14 1446.8075 0.42 ;
      RECT  1447.5075 0.14 1449.6675 0.42 ;
      RECT  1450.3675 0.14 1452.5275 0.42 ;
      RECT  1453.2275 0.14 1455.3875 0.42 ;
      RECT  1456.0875 0.14 1458.2475 0.42 ;
      RECT  1458.9475 0.14 1461.1075 0.42 ;
      RECT  1461.8075 0.14 1463.9675 0.42 ;
      RECT  1464.6675 0.14 1466.8275 0.42 ;
      RECT  1467.5275 0.14 1469.6875 0.42 ;
      RECT  1470.3875 0.14 1472.5475 0.42 ;
      RECT  1473.2475 0.14 1475.4075 0.42 ;
      RECT  1476.1075 0.14 1478.2675 0.42 ;
      RECT  1478.9675 0.14 1481.1275 0.42 ;
      RECT  1481.8275 0.14 1483.9875 0.42 ;
      RECT  1484.6875 0.14 1486.8475 0.42 ;
      RECT  1487.5475 0.14 1489.7075 0.42 ;
      RECT  1490.4075 0.14 1492.5675 0.42 ;
      RECT  1493.2675 0.14 1495.4275 0.42 ;
      RECT  1496.1275 0.14 1498.2875 0.42 ;
      RECT  1498.9875 0.14 1501.1475 0.42 ;
      RECT  1501.8475 0.14 1504.0075 0.42 ;
      RECT  1504.7075 0.14 1506.8675 0.42 ;
      RECT  1507.5675 0.14 1509.7275 0.42 ;
      RECT  1510.4275 0.14 1512.5875 0.42 ;
      RECT  1513.2875 0.14 1515.4475 0.42 ;
      RECT  1516.1475 0.14 1518.3075 0.42 ;
      RECT  1519.0075 0.14 1521.1675 0.42 ;
      RECT  1521.8675 0.14 1524.0275 0.42 ;
      RECT  1524.7275 0.14 1526.8875 0.42 ;
      RECT  1527.5875 0.14 1529.7475 0.42 ;
      RECT  1530.4475 0.14 1532.6075 0.42 ;
      RECT  1533.3075 0.14 1535.4675 0.42 ;
      RECT  1536.1675 0.14 1538.3275 0.42 ;
      RECT  1539.0275 0.14 1541.1875 0.42 ;
      RECT  1541.8875 0.14 1544.0475 0.42 ;
      RECT  1544.7475 0.14 1546.9075 0.42 ;
      RECT  1547.6075 0.14 1549.7675 0.42 ;
      RECT  1550.4675 0.14 1552.6275 0.42 ;
      RECT  1553.3275 0.14 1555.4875 0.42 ;
      RECT  1556.1875 0.14 1558.3475 0.42 ;
      RECT  1559.0475 0.14 1561.2075 0.42 ;
      RECT  1561.9075 0.14 1564.0675 0.42 ;
      RECT  1564.7675 0.14 1566.9275 0.42 ;
      RECT  1567.6275 0.14 1569.7875 0.42 ;
      RECT  1570.4875 0.14 1572.6475 0.42 ;
      RECT  1573.3475 0.14 1575.5075 0.42 ;
      RECT  1576.2075 0.14 1578.3675 0.42 ;
      RECT  1579.0675 0.14 1581.2275 0.42 ;
      RECT  1581.9275 0.14 1584.0875 0.42 ;
      RECT  1584.7875 0.14 1586.9475 0.42 ;
      RECT  1587.6475 0.14 1589.735 0.42 ;
      RECT  0.14 0.42 120.34 171.83 ;
      RECT  120.34 0.42 121.04 171.83 ;
      RECT  121.04 0.42 125.4875 171.83 ;
      RECT  121.04 171.83 125.4875 172.11 ;
      RECT  0.14 171.83 119.2 172.11 ;
      RECT  126.1875 0.42 798.275 171.83 ;
      RECT  798.275 0.42 798.975 171.83 ;
      RECT  798.975 0.42 1589.735 171.83 ;
      RECT  915.6625 171.83 1589.735 172.11 ;
      RECT  799.545 171.83 908.765 172.11 ;
      RECT  909.465 171.83 914.9625 172.11 ;
      RECT  126.1875 171.83 158.1525 172.11 ;
      RECT  158.8525 171.83 159.3275 172.11 ;
      RECT  160.0275 171.83 160.5025 172.11 ;
      RECT  161.2025 171.83 161.6775 172.11 ;
      RECT  162.3775 171.83 162.8525 172.11 ;
      RECT  163.5525 171.83 164.0275 172.11 ;
      RECT  164.7275 171.83 165.2025 172.11 ;
      RECT  165.9025 171.83 166.3775 172.11 ;
      RECT  167.0775 171.83 167.5525 172.11 ;
      RECT  168.2525 171.83 168.7275 172.11 ;
      RECT  169.4275 171.83 169.9025 172.11 ;
      RECT  170.6025 171.83 171.0775 172.11 ;
      RECT  171.7775 171.83 172.2525 172.11 ;
      RECT  172.9525 171.83 173.4275 172.11 ;
      RECT  174.1275 171.83 174.6025 172.11 ;
      RECT  175.3025 171.83 175.7775 172.11 ;
      RECT  176.4775 171.83 176.9525 172.11 ;
      RECT  177.6525 171.83 178.1275 172.11 ;
      RECT  178.8275 171.83 179.3025 172.11 ;
      RECT  180.0025 171.83 180.4775 172.11 ;
      RECT  181.1775 171.83 181.6525 172.11 ;
      RECT  182.3525 171.83 182.8275 172.11 ;
      RECT  183.5275 171.83 184.0025 172.11 ;
      RECT  184.7025 171.83 185.1775 172.11 ;
      RECT  185.8775 171.83 186.3525 172.11 ;
      RECT  187.0525 171.83 187.5275 172.11 ;
      RECT  188.2275 171.83 188.7025 172.11 ;
      RECT  189.4025 171.83 189.8775 172.11 ;
      RECT  190.5775 171.83 191.0525 172.11 ;
      RECT  191.7525 171.83 192.2275 172.11 ;
      RECT  192.9275 171.83 193.4025 172.11 ;
      RECT  194.1025 171.83 194.5775 172.11 ;
      RECT  195.2775 171.83 195.7525 172.11 ;
      RECT  196.4525 171.83 196.9275 172.11 ;
      RECT  197.6275 171.83 198.1025 172.11 ;
      RECT  198.8025 171.83 199.2775 172.11 ;
      RECT  199.9775 171.83 200.4525 172.11 ;
      RECT  201.1525 171.83 201.6275 172.11 ;
      RECT  202.3275 171.83 202.8025 172.11 ;
      RECT  203.5025 171.83 203.9775 172.11 ;
      RECT  204.6775 171.83 205.1525 172.11 ;
      RECT  205.8525 171.83 206.3275 172.11 ;
      RECT  207.0275 171.83 207.5025 172.11 ;
      RECT  208.2025 171.83 208.6775 172.11 ;
      RECT  209.3775 171.83 209.8525 172.11 ;
      RECT  210.5525 171.83 211.0275 172.11 ;
      RECT  211.7275 171.83 212.2025 172.11 ;
      RECT  212.9025 171.83 213.3775 172.11 ;
      RECT  214.0775 171.83 214.5525 172.11 ;
      RECT  215.2525 171.83 215.7275 172.11 ;
      RECT  216.4275 171.83 216.9025 172.11 ;
      RECT  217.6025 171.83 218.0775 172.11 ;
      RECT  218.7775 171.83 219.2525 172.11 ;
      RECT  219.9525 171.83 220.4275 172.11 ;
      RECT  221.1275 171.83 221.6025 172.11 ;
      RECT  222.3025 171.83 222.7775 172.11 ;
      RECT  223.4775 171.83 223.9525 172.11 ;
      RECT  224.6525 171.83 225.1275 172.11 ;
      RECT  225.8275 171.83 226.3025 172.11 ;
      RECT  227.0025 171.83 227.4775 172.11 ;
      RECT  228.1775 171.83 228.6525 172.11 ;
      RECT  229.3525 171.83 229.8275 172.11 ;
      RECT  230.5275 171.83 231.0025 172.11 ;
      RECT  231.7025 171.83 232.1775 172.11 ;
      RECT  232.8775 171.83 233.3525 172.11 ;
      RECT  234.0525 171.83 234.5275 172.11 ;
      RECT  235.2275 171.83 235.7025 172.11 ;
      RECT  236.4025 171.83 236.8775 172.11 ;
      RECT  237.5775 171.83 238.0525 172.11 ;
      RECT  238.7525 171.83 239.2275 172.11 ;
      RECT  239.9275 171.83 240.4025 172.11 ;
      RECT  241.1025 171.83 241.5775 172.11 ;
      RECT  242.2775 171.83 242.7525 172.11 ;
      RECT  243.4525 171.83 243.9275 172.11 ;
      RECT  244.6275 171.83 245.1025 172.11 ;
      RECT  245.8025 171.83 246.2775 172.11 ;
      RECT  246.9775 171.83 247.4525 172.11 ;
      RECT  248.1525 171.83 248.6275 172.11 ;
      RECT  249.3275 171.83 249.8025 172.11 ;
      RECT  250.5025 171.83 250.9775 172.11 ;
      RECT  251.6775 171.83 252.1525 172.11 ;
      RECT  252.8525 171.83 253.3275 172.11 ;
      RECT  254.0275 171.83 254.5025 172.11 ;
      RECT  255.2025 171.83 255.6775 172.11 ;
      RECT  256.3775 171.83 256.8525 172.11 ;
      RECT  257.5525 171.83 258.0275 172.11 ;
      RECT  258.7275 171.83 259.2025 172.11 ;
      RECT  259.9025 171.83 260.3775 172.11 ;
      RECT  261.0775 171.83 261.5525 172.11 ;
      RECT  262.2525 171.83 262.7275 172.11 ;
      RECT  263.4275 171.83 263.9025 172.11 ;
      RECT  264.6025 171.83 265.0775 172.11 ;
      RECT  265.7775 171.83 266.2525 172.11 ;
      RECT  266.9525 171.83 267.4275 172.11 ;
      RECT  268.1275 171.83 268.6025 172.11 ;
      RECT  269.3025 171.83 269.7775 172.11 ;
      RECT  270.4775 171.83 270.9525 172.11 ;
      RECT  271.6525 171.83 272.1275 172.11 ;
      RECT  272.8275 171.83 273.3025 172.11 ;
      RECT  274.0025 171.83 274.4775 172.11 ;
      RECT  275.1775 171.83 275.6525 172.11 ;
      RECT  276.3525 171.83 276.8275 172.11 ;
      RECT  277.5275 171.83 278.0025 172.11 ;
      RECT  278.7025 171.83 279.1775 172.11 ;
      RECT  279.8775 171.83 280.3525 172.11 ;
      RECT  281.0525 171.83 281.5275 172.11 ;
      RECT  282.2275 171.83 282.7025 172.11 ;
      RECT  283.4025 171.83 283.8775 172.11 ;
      RECT  284.5775 171.83 285.0525 172.11 ;
      RECT  285.7525 171.83 286.2275 172.11 ;
      RECT  286.9275 171.83 287.4025 172.11 ;
      RECT  288.1025 171.83 288.5775 172.11 ;
      RECT  289.2775 171.83 289.7525 172.11 ;
      RECT  290.4525 171.83 290.9275 172.11 ;
      RECT  291.6275 171.83 292.1025 172.11 ;
      RECT  292.8025 171.83 293.2775 172.11 ;
      RECT  293.9775 171.83 294.4525 172.11 ;
      RECT  295.1525 171.83 295.6275 172.11 ;
      RECT  296.3275 171.83 296.8025 172.11 ;
      RECT  297.5025 171.83 297.9775 172.11 ;
      RECT  298.6775 171.83 299.1525 172.11 ;
      RECT  299.8525 171.83 300.3275 172.11 ;
      RECT  301.0275 171.83 301.5025 172.11 ;
      RECT  302.2025 171.83 302.6775 172.11 ;
      RECT  303.3775 171.83 303.8525 172.11 ;
      RECT  304.5525 171.83 305.0275 172.11 ;
      RECT  305.7275 171.83 306.2025 172.11 ;
      RECT  306.9025 171.83 307.3775 172.11 ;
      RECT  308.0775 171.83 308.5525 172.11 ;
      RECT  309.2525 171.83 309.7275 172.11 ;
      RECT  310.4275 171.83 310.9025 172.11 ;
      RECT  311.6025 171.83 312.0775 172.11 ;
      RECT  312.7775 171.83 313.2525 172.11 ;
      RECT  313.9525 171.83 314.4275 172.11 ;
      RECT  315.1275 171.83 315.6025 172.11 ;
      RECT  316.3025 171.83 316.7775 172.11 ;
      RECT  317.4775 171.83 317.9525 172.11 ;
      RECT  318.6525 171.83 319.1275 172.11 ;
      RECT  319.8275 171.83 320.3025 172.11 ;
      RECT  321.0025 171.83 321.4775 172.11 ;
      RECT  322.1775 171.83 322.6525 172.11 ;
      RECT  323.3525 171.83 323.8275 172.11 ;
      RECT  324.5275 171.83 325.0025 172.11 ;
      RECT  325.7025 171.83 326.1775 172.11 ;
      RECT  326.8775 171.83 327.3525 172.11 ;
      RECT  328.0525 171.83 328.5275 172.11 ;
      RECT  329.2275 171.83 329.7025 172.11 ;
      RECT  330.4025 171.83 330.8775 172.11 ;
      RECT  331.5775 171.83 332.0525 172.11 ;
      RECT  332.7525 171.83 333.2275 172.11 ;
      RECT  333.9275 171.83 334.4025 172.11 ;
      RECT  335.1025 171.83 335.5775 172.11 ;
      RECT  336.2775 171.83 336.7525 172.11 ;
      RECT  337.4525 171.83 337.9275 172.11 ;
      RECT  338.6275 171.83 339.1025 172.11 ;
      RECT  339.8025 171.83 340.2775 172.11 ;
      RECT  340.9775 171.83 341.4525 172.11 ;
      RECT  342.1525 171.83 342.6275 172.11 ;
      RECT  343.3275 171.83 343.8025 172.11 ;
      RECT  344.5025 171.83 344.9775 172.11 ;
      RECT  345.6775 171.83 346.1525 172.11 ;
      RECT  346.8525 171.83 347.3275 172.11 ;
      RECT  348.0275 171.83 348.5025 172.11 ;
      RECT  349.2025 171.83 349.6775 172.11 ;
      RECT  350.3775 171.83 350.8525 172.11 ;
      RECT  351.5525 171.83 352.0275 172.11 ;
      RECT  352.7275 171.83 353.2025 172.11 ;
      RECT  353.9025 171.83 354.3775 172.11 ;
      RECT  355.0775 171.83 355.5525 172.11 ;
      RECT  356.2525 171.83 356.7275 172.11 ;
      RECT  357.4275 171.83 357.9025 172.11 ;
      RECT  358.6025 171.83 359.0775 172.11 ;
      RECT  359.7775 171.83 360.2525 172.11 ;
      RECT  360.9525 171.83 361.4275 172.11 ;
      RECT  362.1275 171.83 362.6025 172.11 ;
      RECT  363.3025 171.83 363.7775 172.11 ;
      RECT  364.4775 171.83 364.9525 172.11 ;
      RECT  365.6525 171.83 366.1275 172.11 ;
      RECT  366.8275 171.83 367.3025 172.11 ;
      RECT  368.0025 171.83 368.4775 172.11 ;
      RECT  369.1775 171.83 369.6525 172.11 ;
      RECT  370.3525 171.83 370.8275 172.11 ;
      RECT  371.5275 171.83 372.0025 172.11 ;
      RECT  372.7025 171.83 373.1775 172.11 ;
      RECT  373.8775 171.83 374.3525 172.11 ;
      RECT  375.0525 171.83 375.5275 172.11 ;
      RECT  376.2275 171.83 376.7025 172.11 ;
      RECT  377.4025 171.83 377.8775 172.11 ;
      RECT  378.5775 171.83 379.0525 172.11 ;
      RECT  379.7525 171.83 380.2275 172.11 ;
      RECT  380.9275 171.83 381.4025 172.11 ;
      RECT  382.1025 171.83 382.5775 172.11 ;
      RECT  383.2775 171.83 383.7525 172.11 ;
      RECT  384.4525 171.83 384.9275 172.11 ;
      RECT  385.6275 171.83 386.1025 172.11 ;
      RECT  386.8025 171.83 387.2775 172.11 ;
      RECT  387.9775 171.83 388.4525 172.11 ;
      RECT  389.1525 171.83 389.6275 172.11 ;
      RECT  390.3275 171.83 390.8025 172.11 ;
      RECT  391.5025 171.83 391.9775 172.11 ;
      RECT  392.6775 171.83 393.1525 172.11 ;
      RECT  393.8525 171.83 394.3275 172.11 ;
      RECT  395.0275 171.83 395.5025 172.11 ;
      RECT  396.2025 171.83 396.6775 172.11 ;
      RECT  397.3775 171.83 397.8525 172.11 ;
      RECT  398.5525 171.83 399.0275 172.11 ;
      RECT  399.7275 171.83 400.2025 172.11 ;
      RECT  400.9025 171.83 401.3775 172.11 ;
      RECT  402.0775 171.83 402.5525 172.11 ;
      RECT  403.2525 171.83 403.7275 172.11 ;
      RECT  404.4275 171.83 404.9025 172.11 ;
      RECT  405.6025 171.83 406.0775 172.11 ;
      RECT  406.7775 171.83 407.2525 172.11 ;
      RECT  407.9525 171.83 408.4275 172.11 ;
      RECT  409.1275 171.83 409.6025 172.11 ;
      RECT  410.3025 171.83 410.7775 172.11 ;
      RECT  411.4775 171.83 411.9525 172.11 ;
      RECT  412.6525 171.83 413.1275 172.11 ;
      RECT  413.8275 171.83 414.3025 172.11 ;
      RECT  415.0025 171.83 415.4775 172.11 ;
      RECT  416.1775 171.83 416.6525 172.11 ;
      RECT  417.3525 171.83 417.8275 172.11 ;
      RECT  418.5275 171.83 419.0025 172.11 ;
      RECT  419.7025 171.83 420.1775 172.11 ;
      RECT  420.8775 171.83 421.3525 172.11 ;
      RECT  422.0525 171.83 422.5275 172.11 ;
      RECT  423.2275 171.83 423.7025 172.11 ;
      RECT  424.4025 171.83 424.8775 172.11 ;
      RECT  425.5775 171.83 426.0525 172.11 ;
      RECT  426.7525 171.83 427.2275 172.11 ;
      RECT  427.9275 171.83 428.4025 172.11 ;
      RECT  429.1025 171.83 429.5775 172.11 ;
      RECT  430.2775 171.83 430.7525 172.11 ;
      RECT  431.4525 171.83 431.9275 172.11 ;
      RECT  432.6275 171.83 433.1025 172.11 ;
      RECT  433.8025 171.83 434.2775 172.11 ;
      RECT  434.9775 171.83 435.4525 172.11 ;
      RECT  436.1525 171.83 436.6275 172.11 ;
      RECT  437.3275 171.83 437.8025 172.11 ;
      RECT  438.5025 171.83 438.9775 172.11 ;
      RECT  439.6775 171.83 440.1525 172.11 ;
      RECT  440.8525 171.83 441.3275 172.11 ;
      RECT  442.0275 171.83 442.5025 172.11 ;
      RECT  443.2025 171.83 443.6775 172.11 ;
      RECT  444.3775 171.83 444.8525 172.11 ;
      RECT  445.5525 171.83 446.0275 172.11 ;
      RECT  446.7275 171.83 447.2025 172.11 ;
      RECT  447.9025 171.83 448.3775 172.11 ;
      RECT  449.0775 171.83 449.5525 172.11 ;
      RECT  450.2525 171.83 450.7275 172.11 ;
      RECT  451.4275 171.83 451.9025 172.11 ;
      RECT  452.6025 171.83 453.0775 172.11 ;
      RECT  453.7775 171.83 454.2525 172.11 ;
      RECT  454.9525 171.83 455.4275 172.11 ;
      RECT  456.1275 171.83 456.6025 172.11 ;
      RECT  457.3025 171.83 457.7775 172.11 ;
      RECT  458.4775 171.83 458.9525 172.11 ;
      RECT  459.6525 171.83 460.1275 172.11 ;
      RECT  460.8275 171.83 461.3025 172.11 ;
      RECT  462.0025 171.83 462.4775 172.11 ;
      RECT  463.1775 171.83 463.6525 172.11 ;
      RECT  464.3525 171.83 464.8275 172.11 ;
      RECT  465.5275 171.83 466.0025 172.11 ;
      RECT  466.7025 171.83 467.1775 172.11 ;
      RECT  467.8775 171.83 468.3525 172.11 ;
      RECT  469.0525 171.83 469.5275 172.11 ;
      RECT  470.2275 171.83 470.7025 172.11 ;
      RECT  471.4025 171.83 471.8775 172.11 ;
      RECT  472.5775 171.83 473.0525 172.11 ;
      RECT  473.7525 171.83 474.2275 172.11 ;
      RECT  474.9275 171.83 475.4025 172.11 ;
      RECT  476.1025 171.83 476.5775 172.11 ;
      RECT  477.2775 171.83 477.7525 172.11 ;
      RECT  478.4525 171.83 478.9275 172.11 ;
      RECT  479.6275 171.83 480.1025 172.11 ;
      RECT  480.8025 171.83 481.2775 172.11 ;
      RECT  481.9775 171.83 482.4525 172.11 ;
      RECT  483.1525 171.83 483.6275 172.11 ;
      RECT  484.3275 171.83 484.8025 172.11 ;
      RECT  485.5025 171.83 485.9775 172.11 ;
      RECT  486.6775 171.83 487.1525 172.11 ;
      RECT  487.8525 171.83 488.3275 172.11 ;
      RECT  489.0275 171.83 489.5025 172.11 ;
      RECT  490.2025 171.83 490.6775 172.11 ;
      RECT  491.3775 171.83 491.8525 172.11 ;
      RECT  492.5525 171.83 493.0275 172.11 ;
      RECT  493.7275 171.83 494.2025 172.11 ;
      RECT  494.9025 171.83 495.3775 172.11 ;
      RECT  496.0775 171.83 496.5525 172.11 ;
      RECT  497.2525 171.83 497.7275 172.11 ;
      RECT  498.4275 171.83 498.9025 172.11 ;
      RECT  499.6025 171.83 500.0775 172.11 ;
      RECT  500.7775 171.83 501.2525 172.11 ;
      RECT  501.9525 171.83 502.4275 172.11 ;
      RECT  503.1275 171.83 503.6025 172.11 ;
      RECT  504.3025 171.83 504.7775 172.11 ;
      RECT  505.4775 171.83 505.9525 172.11 ;
      RECT  506.6525 171.83 507.1275 172.11 ;
      RECT  507.8275 171.83 508.3025 172.11 ;
      RECT  509.0025 171.83 509.4775 172.11 ;
      RECT  510.1775 171.83 510.6525 172.11 ;
      RECT  511.3525 171.83 511.8275 172.11 ;
      RECT  512.5275 171.83 513.0025 172.11 ;
      RECT  513.7025 171.83 514.1775 172.11 ;
      RECT  514.8775 171.83 515.3525 172.11 ;
      RECT  516.0525 171.83 516.5275 172.11 ;
      RECT  517.2275 171.83 517.7025 172.11 ;
      RECT  518.4025 171.83 518.8775 172.11 ;
      RECT  519.5775 171.83 520.0525 172.11 ;
      RECT  520.7525 171.83 521.2275 172.11 ;
      RECT  521.9275 171.83 522.4025 172.11 ;
      RECT  523.1025 171.83 523.5775 172.11 ;
      RECT  524.2775 171.83 524.7525 172.11 ;
      RECT  525.4525 171.83 525.9275 172.11 ;
      RECT  526.6275 171.83 527.1025 172.11 ;
      RECT  527.8025 171.83 528.2775 172.11 ;
      RECT  528.9775 171.83 529.4525 172.11 ;
      RECT  530.1525 171.83 530.6275 172.11 ;
      RECT  531.3275 171.83 531.8025 172.11 ;
      RECT  532.5025 171.83 532.9775 172.11 ;
      RECT  533.6775 171.83 534.1525 172.11 ;
      RECT  534.8525 171.83 535.3275 172.11 ;
      RECT  536.0275 171.83 536.5025 172.11 ;
      RECT  537.2025 171.83 537.6775 172.11 ;
      RECT  538.3775 171.83 538.8525 172.11 ;
      RECT  539.5525 171.83 540.0275 172.11 ;
      RECT  540.7275 171.83 541.2025 172.11 ;
      RECT  541.9025 171.83 542.3775 172.11 ;
      RECT  543.0775 171.83 543.5525 172.11 ;
      RECT  544.2525 171.83 544.7275 172.11 ;
      RECT  545.4275 171.83 545.9025 172.11 ;
      RECT  546.6025 171.83 547.0775 172.11 ;
      RECT  547.7775 171.83 548.2525 172.11 ;
      RECT  548.9525 171.83 549.4275 172.11 ;
      RECT  550.1275 171.83 550.6025 172.11 ;
      RECT  551.3025 171.83 551.7775 172.11 ;
      RECT  552.4775 171.83 552.9525 172.11 ;
      RECT  553.6525 171.83 554.1275 172.11 ;
      RECT  554.8275 171.83 555.3025 172.11 ;
      RECT  556.0025 171.83 556.4775 172.11 ;
      RECT  557.1775 171.83 557.6525 172.11 ;
      RECT  558.3525 171.83 558.8275 172.11 ;
      RECT  559.5275 171.83 560.0025 172.11 ;
      RECT  560.7025 171.83 561.1775 172.11 ;
      RECT  561.8775 171.83 562.3525 172.11 ;
      RECT  563.0525 171.83 563.5275 172.11 ;
      RECT  564.2275 171.83 564.7025 172.11 ;
      RECT  565.4025 171.83 565.8775 172.11 ;
      RECT  566.5775 171.83 567.0525 172.11 ;
      RECT  567.7525 171.83 568.2275 172.11 ;
      RECT  568.9275 171.83 569.4025 172.11 ;
      RECT  570.1025 171.83 570.5775 172.11 ;
      RECT  571.2775 171.83 571.7525 172.11 ;
      RECT  572.4525 171.83 572.9275 172.11 ;
      RECT  573.6275 171.83 574.1025 172.11 ;
      RECT  574.8025 171.83 575.2775 172.11 ;
      RECT  575.9775 171.83 576.4525 172.11 ;
      RECT  577.1525 171.83 577.6275 172.11 ;
      RECT  578.3275 171.83 578.8025 172.11 ;
      RECT  579.5025 171.83 579.9775 172.11 ;
      RECT  580.6775 171.83 581.1525 172.11 ;
      RECT  581.8525 171.83 582.3275 172.11 ;
      RECT  583.0275 171.83 583.5025 172.11 ;
      RECT  584.2025 171.83 584.6775 172.11 ;
      RECT  585.3775 171.83 585.8525 172.11 ;
      RECT  586.5525 171.83 587.0275 172.11 ;
      RECT  587.7275 171.83 588.2025 172.11 ;
      RECT  588.9025 171.83 589.3775 172.11 ;
      RECT  590.0775 171.83 590.5525 172.11 ;
      RECT  591.2525 171.83 591.7275 172.11 ;
      RECT  592.4275 171.83 592.9025 172.11 ;
      RECT  593.6025 171.83 594.0775 172.11 ;
      RECT  594.7775 171.83 595.2525 172.11 ;
      RECT  595.9525 171.83 596.4275 172.11 ;
      RECT  597.1275 171.83 597.6025 172.11 ;
      RECT  598.3025 171.83 598.7775 172.11 ;
      RECT  599.4775 171.83 599.9525 172.11 ;
      RECT  600.6525 171.83 601.1275 172.11 ;
      RECT  601.8275 171.83 602.3025 172.11 ;
      RECT  603.0025 171.83 603.4775 172.11 ;
      RECT  604.1775 171.83 604.6525 172.11 ;
      RECT  605.3525 171.83 605.8275 172.11 ;
      RECT  606.5275 171.83 607.0025 172.11 ;
      RECT  607.7025 171.83 608.1775 172.11 ;
      RECT  608.8775 171.83 609.3525 172.11 ;
      RECT  610.0525 171.83 610.5275 172.11 ;
      RECT  611.2275 171.83 611.7025 172.11 ;
      RECT  612.4025 171.83 612.8775 172.11 ;
      RECT  613.5775 171.83 614.0525 172.11 ;
      RECT  614.7525 171.83 615.2275 172.11 ;
      RECT  615.9275 171.83 616.4025 172.11 ;
      RECT  617.1025 171.83 617.5775 172.11 ;
      RECT  618.2775 171.83 618.7525 172.11 ;
      RECT  619.4525 171.83 619.9275 172.11 ;
      RECT  620.6275 171.83 621.1025 172.11 ;
      RECT  621.8025 171.83 622.2775 172.11 ;
      RECT  622.9775 171.83 623.4525 172.11 ;
      RECT  624.1525 171.83 624.6275 172.11 ;
      RECT  625.3275 171.83 625.8025 172.11 ;
      RECT  626.5025 171.83 626.9775 172.11 ;
      RECT  627.6775 171.83 628.1525 172.11 ;
      RECT  628.8525 171.83 629.3275 172.11 ;
      RECT  630.0275 171.83 630.5025 172.11 ;
      RECT  631.2025 171.83 631.6775 172.11 ;
      RECT  632.3775 171.83 632.8525 172.11 ;
      RECT  633.5525 171.83 634.0275 172.11 ;
      RECT  634.7275 171.83 635.2025 172.11 ;
      RECT  635.9025 171.83 636.3775 172.11 ;
      RECT  637.0775 171.83 637.5525 172.11 ;
      RECT  638.2525 171.83 638.7275 172.11 ;
      RECT  639.4275 171.83 639.9025 172.11 ;
      RECT  640.6025 171.83 641.0775 172.11 ;
      RECT  641.7775 171.83 642.2525 172.11 ;
      RECT  642.9525 171.83 643.4275 172.11 ;
      RECT  644.1275 171.83 644.6025 172.11 ;
      RECT  645.3025 171.83 645.7775 172.11 ;
      RECT  646.4775 171.83 646.9525 172.11 ;
      RECT  647.6525 171.83 648.1275 172.11 ;
      RECT  648.8275 171.83 649.3025 172.11 ;
      RECT  650.0025 171.83 650.4775 172.11 ;
      RECT  651.1775 171.83 651.6525 172.11 ;
      RECT  652.3525 171.83 652.8275 172.11 ;
      RECT  653.5275 171.83 654.0025 172.11 ;
      RECT  654.7025 171.83 655.1775 172.11 ;
      RECT  655.8775 171.83 656.3525 172.11 ;
      RECT  657.0525 171.83 657.5275 172.11 ;
      RECT  658.2275 171.83 658.7025 172.11 ;
      RECT  659.4025 171.83 659.8775 172.11 ;
      RECT  660.5775 171.83 661.0525 172.11 ;
      RECT  661.7525 171.83 662.2275 172.11 ;
      RECT  662.9275 171.83 663.4025 172.11 ;
      RECT  664.1025 171.83 664.5775 172.11 ;
      RECT  665.2775 171.83 665.7525 172.11 ;
      RECT  666.4525 171.83 666.9275 172.11 ;
      RECT  667.6275 171.83 668.1025 172.11 ;
      RECT  668.8025 171.83 669.2775 172.11 ;
      RECT  669.9775 171.83 670.4525 172.11 ;
      RECT  671.1525 171.83 671.6275 172.11 ;
      RECT  672.3275 171.83 672.8025 172.11 ;
      RECT  673.5025 171.83 673.9775 172.11 ;
      RECT  674.6775 171.83 675.1525 172.11 ;
      RECT  675.8525 171.83 676.3275 172.11 ;
      RECT  677.0275 171.83 677.5025 172.11 ;
      RECT  678.2025 171.83 678.6775 172.11 ;
      RECT  679.3775 171.83 679.8525 172.11 ;
      RECT  680.5525 171.83 681.0275 172.11 ;
      RECT  681.7275 171.83 682.2025 172.11 ;
      RECT  682.9025 171.83 683.3775 172.11 ;
      RECT  684.0775 171.83 684.5525 172.11 ;
      RECT  685.2525 171.83 685.7275 172.11 ;
      RECT  686.4275 171.83 686.9025 172.11 ;
      RECT  687.6025 171.83 688.0775 172.11 ;
      RECT  688.7775 171.83 689.2525 172.11 ;
      RECT  689.9525 171.83 690.4275 172.11 ;
      RECT  691.1275 171.83 691.6025 172.11 ;
      RECT  692.3025 171.83 692.7775 172.11 ;
      RECT  693.4775 171.83 693.9525 172.11 ;
      RECT  694.6525 171.83 695.1275 172.11 ;
      RECT  695.8275 171.83 696.3025 172.11 ;
      RECT  697.0025 171.83 697.4775 172.11 ;
      RECT  698.1775 171.83 698.6525 172.11 ;
      RECT  699.3525 171.83 699.8275 172.11 ;
      RECT  700.5275 171.83 701.0025 172.11 ;
      RECT  701.7025 171.83 702.1775 172.11 ;
      RECT  702.8775 171.83 703.3525 172.11 ;
      RECT  704.0525 171.83 704.5275 172.11 ;
      RECT  705.2275 171.83 705.7025 172.11 ;
      RECT  706.4025 171.83 706.8775 172.11 ;
      RECT  707.5775 171.83 708.0525 172.11 ;
      RECT  708.7525 171.83 709.2275 172.11 ;
      RECT  709.9275 171.83 710.4025 172.11 ;
      RECT  711.1025 171.83 711.5775 172.11 ;
      RECT  712.2775 171.83 712.7525 172.11 ;
      RECT  713.4525 171.83 713.9275 172.11 ;
      RECT  714.6275 171.83 715.1025 172.11 ;
      RECT  715.8025 171.83 716.2775 172.11 ;
      RECT  716.9775 171.83 717.4525 172.11 ;
      RECT  718.1525 171.83 718.6275 172.11 ;
      RECT  719.3275 171.83 719.8025 172.11 ;
      RECT  720.5025 171.83 720.9775 172.11 ;
      RECT  721.6775 171.83 722.1525 172.11 ;
      RECT  722.8525 171.83 723.3275 172.11 ;
      RECT  724.0275 171.83 724.5025 172.11 ;
      RECT  725.2025 171.83 725.6775 172.11 ;
      RECT  726.3775 171.83 726.8525 172.11 ;
      RECT  727.5525 171.83 728.0275 172.11 ;
      RECT  728.7275 171.83 729.2025 172.11 ;
      RECT  729.9025 171.83 730.3775 172.11 ;
      RECT  731.0775 171.83 731.5525 172.11 ;
      RECT  732.2525 171.83 732.7275 172.11 ;
      RECT  733.4275 171.83 733.9025 172.11 ;
      RECT  734.6025 171.83 735.0775 172.11 ;
      RECT  735.7775 171.83 736.2525 172.11 ;
      RECT  736.9525 171.83 737.4275 172.11 ;
      RECT  738.1275 171.83 738.6025 172.11 ;
      RECT  739.3025 171.83 739.7775 172.11 ;
      RECT  740.4775 171.83 740.9525 172.11 ;
      RECT  741.6525 171.83 742.1275 172.11 ;
      RECT  742.8275 171.83 743.3025 172.11 ;
      RECT  744.0025 171.83 744.4775 172.11 ;
      RECT  745.1775 171.83 745.6525 172.11 ;
      RECT  746.3525 171.83 746.8275 172.11 ;
      RECT  747.5275 171.83 748.0025 172.11 ;
      RECT  748.7025 171.83 749.1775 172.11 ;
      RECT  749.8775 171.83 750.3525 172.11 ;
      RECT  751.0525 171.83 751.5275 172.11 ;
      RECT  752.2275 171.83 752.7025 172.11 ;
      RECT  753.4025 171.83 753.8775 172.11 ;
      RECT  754.5775 171.83 755.0525 172.11 ;
      RECT  755.7525 171.83 756.2275 172.11 ;
      RECT  756.9275 171.83 757.4025 172.11 ;
      RECT  758.1025 171.83 758.5775 172.11 ;
      RECT  759.2775 171.83 797.99 172.11 ;
   END
END    sram_0rw1r1w_512_16_freepdk45
END    LIBRARY
