VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_1rw0r0w_32_128_freepdk45
   CLASS BLOCK ;
   SIZE 119.29 BY 117.815 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  27.9825 0.0 28.1225 0.14 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  30.8425 0.0 30.9825 0.14 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  33.7025 0.0 33.8425 0.14 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  36.5625 0.0 36.7025 0.14 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  39.4225 0.0 39.5625 0.14 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  42.2825 0.0 42.4225 0.14 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  45.1425 0.0 45.2825 0.14 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  48.0025 0.0 48.1425 0.14 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  50.8625 0.0 51.0025 0.14 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  53.7225 0.0 53.8625 0.14 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  56.5825 0.0 56.7225 0.14 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  59.4425 0.0 59.5825 0.14 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  62.3025 0.0 62.4425 0.14 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  65.1625 0.0 65.3025 0.14 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  68.0225 0.0 68.1625 0.14 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  70.8825 0.0 71.0225 0.14 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  73.7425 0.0 73.8825 0.14 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  76.6025 0.0 76.7425 0.14 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  79.4625 0.0 79.6025 0.14 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  82.3225 0.0 82.4625 0.14 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  85.1825 0.0 85.3225 0.14 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  88.0425 0.0 88.1825 0.14 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  90.9025 0.0 91.0425 0.14 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  93.7625 0.0 93.9025 0.14 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  96.6225 0.0 96.7625 0.14 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  99.4825 0.0 99.6225 0.14 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  102.3425 0.0 102.4825 0.14 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  105.2025 0.0 105.3425 0.14 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  108.0625 0.0 108.2025 0.14 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  110.9225 0.0 111.0625 0.14 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  113.7825 0.0 113.9225 0.14 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  116.6425 0.0 116.7825 0.14 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  25.1225 0.0 25.2625 0.14 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 51.7 0.14 51.84 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 54.43 0.14 54.57 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 56.64 0.14 56.78 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 59.37 0.14 59.51 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 61.58 0.14 61.72 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 64.31 0.14 64.45 ;
      END
   END addr0[6]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 6.98 0.14 7.12 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 9.71 0.14 9.85 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  9.84 0.0 9.98 0.14 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  39.905 0.0 40.045 0.14 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  40.7425 0.0 40.8825 0.14 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  42.725 0.0 42.865 0.14 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  43.5625 0.0 43.7025 0.14 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  45.545 0.0 45.685 0.14 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  46.3825 0.0 46.5225 0.14 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  47.245 0.0 47.385 0.14 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  49.2025 0.0 49.3425 0.14 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  50.105 0.0 50.245 0.14 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  52.0225 0.0 52.1625 0.14 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  52.965 0.0 53.105 0.14 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  54.8425 0.0 54.9825 0.14 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  55.825 0.0 55.965 0.14 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  57.6625 0.0 57.8025 0.14 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  58.685 0.0 58.825 0.14 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  60.4825 0.0 60.6225 0.14 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  61.545 0.0 61.685 0.14 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  63.3025 0.0 63.4425 0.14 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  64.405 0.0 64.545 0.14 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  66.1225 0.0 66.2625 0.14 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  67.265 0.0 67.405 0.14 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  68.9425 0.0 69.0825 0.14 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  70.1175 0.0 70.2575 0.14 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  71.7625 0.0 71.9025 0.14 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  72.9375 0.0 73.0775 0.14 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  74.5825 0.0 74.7225 0.14 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  75.7575 0.0 75.8975 0.14 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  77.4025 0.0 77.5425 0.14 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  78.705 0.0 78.845 0.14 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  80.2225 0.0 80.3625 0.14 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  81.565 0.0 81.705 0.14 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  83.0425 0.0 83.1825 0.14 ;
      END
   END dout0[31]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 119.15 117.675 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 119.15 117.675 ;
   LAYER  metal3 ;
      RECT  0.28 0.14 119.15 51.56 ;
      RECT  0.28 51.56 119.15 51.98 ;
      RECT  0.28 51.98 119.15 117.675 ;
      RECT  0.14 51.98 0.28 54.29 ;
      RECT  0.14 54.71 0.28 56.5 ;
      RECT  0.14 56.92 0.28 59.23 ;
      RECT  0.14 59.65 0.28 61.44 ;
      RECT  0.14 61.86 0.28 64.17 ;
      RECT  0.14 64.59 0.28 117.675 ;
      RECT  0.14 0.14 0.28 6.84 ;
      RECT  0.14 7.26 0.28 9.57 ;
      RECT  0.14 9.99 0.28 51.56 ;
   LAYER  metal4 ;
      RECT  0.14 0.42 27.7025 117.675 ;
      RECT  27.7025 0.42 28.4025 117.675 ;
      RECT  28.4025 0.42 119.15 117.675 ;
      RECT  28.4025 0.14 30.5625 0.42 ;
      RECT  31.2625 0.14 33.4225 0.42 ;
      RECT  34.1225 0.14 36.2825 0.42 ;
      RECT  36.9825 0.14 39.1425 0.42 ;
      RECT  85.6025 0.14 87.7625 0.42 ;
      RECT  88.4625 0.14 90.6225 0.42 ;
      RECT  91.3225 0.14 93.4825 0.42 ;
      RECT  94.1825 0.14 96.3425 0.42 ;
      RECT  97.0425 0.14 99.2025 0.42 ;
      RECT  99.9025 0.14 102.0625 0.42 ;
      RECT  102.7625 0.14 104.9225 0.42 ;
      RECT  105.6225 0.14 107.7825 0.42 ;
      RECT  108.4825 0.14 110.6425 0.42 ;
      RECT  111.3425 0.14 113.5025 0.42 ;
      RECT  114.2025 0.14 116.3625 0.42 ;
      RECT  117.0625 0.14 119.15 0.42 ;
      RECT  25.5425 0.14 27.7025 0.42 ;
      RECT  0.14 0.14 9.56 0.42 ;
      RECT  10.26 0.14 24.8425 0.42 ;
      RECT  40.325 0.14 40.4625 0.42 ;
      RECT  41.1625 0.14 42.0025 0.42 ;
      RECT  43.145 0.14 43.2825 0.42 ;
      RECT  43.9825 0.14 44.8625 0.42 ;
      RECT  45.965 0.14 46.1025 0.42 ;
      RECT  46.8025 0.14 46.965 0.42 ;
      RECT  47.665 0.14 47.7225 0.42 ;
      RECT  48.4225 0.14 48.9225 0.42 ;
      RECT  49.6225 0.14 49.825 0.42 ;
      RECT  50.525 0.14 50.5825 0.42 ;
      RECT  51.2825 0.14 51.7425 0.42 ;
      RECT  52.4425 0.14 52.685 0.42 ;
      RECT  53.385 0.14 53.4425 0.42 ;
      RECT  54.1425 0.14 54.5625 0.42 ;
      RECT  55.2625 0.14 55.545 0.42 ;
      RECT  56.245 0.14 56.3025 0.42 ;
      RECT  57.0025 0.14 57.3825 0.42 ;
      RECT  58.0825 0.14 58.405 0.42 ;
      RECT  59.105 0.14 59.1625 0.42 ;
      RECT  59.8625 0.14 60.2025 0.42 ;
      RECT  60.9025 0.14 61.265 0.42 ;
      RECT  61.965 0.14 62.0225 0.42 ;
      RECT  62.7225 0.14 63.0225 0.42 ;
      RECT  63.7225 0.14 64.125 0.42 ;
      RECT  64.825 0.14 64.8825 0.42 ;
      RECT  65.5825 0.14 65.8425 0.42 ;
      RECT  66.5425 0.14 66.985 0.42 ;
      RECT  67.685 0.14 67.7425 0.42 ;
      RECT  68.4425 0.14 68.6625 0.42 ;
      RECT  69.3625 0.14 69.8375 0.42 ;
      RECT  70.5375 0.14 70.6025 0.42 ;
      RECT  71.3025 0.14 71.4825 0.42 ;
      RECT  72.1825 0.14 72.6575 0.42 ;
      RECT  73.3575 0.14 73.4625 0.42 ;
      RECT  74.1625 0.14 74.3025 0.42 ;
      RECT  75.0025 0.14 75.4775 0.42 ;
      RECT  76.1775 0.14 76.3225 0.42 ;
      RECT  77.0225 0.14 77.1225 0.42 ;
      RECT  77.8225 0.14 78.425 0.42 ;
      RECT  79.125 0.14 79.1825 0.42 ;
      RECT  79.8825 0.14 79.9425 0.42 ;
      RECT  80.6425 0.14 81.285 0.42 ;
      RECT  81.985 0.14 82.0425 0.42 ;
      RECT  82.7425 0.14 82.7625 0.42 ;
      RECT  83.4625 0.14 84.9025 0.42 ;
   END
END    sram_1rw0r0w_32_128_freepdk45
END    LIBRARY
