
* cell example_config_freepdk45
* pin csb0
* pin web0
* pin addr0[3]
* pin clk0
* pin dout0[1]
* pin dout0[0]
* pin addr0[2]
* pin addr0[1]
* pin addr0[0]
* pin din0[0]
* pin din0[1]
* pin NWELL
* pin BULK,PWELL
.SUBCKT example_config_freepdk45 7 8 9 10 11 12 13 14 15 16 17 22 23
* net 7 csb0
* net 8 web0
* net 9 addr0[3]
* net 10 clk0
* net 11 dout0[1]
* net 12 dout0[0]
* net 13 addr0[2]
* net 14 addr0[1]
* net 15 addr0[0]
* net 16 din0[0]
* net 17 din0[1]
* net 22 NWELL
* net 23 BULK,PWELL
* cell instance $1 r0 *1 3.15,3.215
X$1 7 1 10 8 2 3 4 6 5 22 23 example_config_freepdk45_control_logic_rw
* cell instance $2 r0 *1 10.94,39.745
X$2 15 18 14 19 13 20 9 21 1 22 23 example_config_freepdk45_row_addr_dff
* cell instance $3 r0 *1 16.66,3.215
X$3 16 25 17 24 1 22 23 example_config_freepdk45_data_dff
* cell instance $7 r0 *1 14.08,10.075
X$7 25 24 3 4 2 12 11 6 5 18 19 20 21 22 23 example_config_freepdk45_bank
.ENDS example_config_freepdk45

* cell example_config_freepdk45_data_dff
* pin din_0
* pin dout_0
* pin din_1
* pin dout_1
* pin clk
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_data_dff 1 2 3 4 5 6 7
* net 1 din_0
* net 2 dout_0
* net 3 din_1
* net 4 dout_1
* net 5 clk
* net 6 vdd
* net 7 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 5 6 7 dff
* cell instance $2 r0 *1 2.86,0
X$2 4 3 5 6 7 dff
.ENDS example_config_freepdk45_data_dff

* cell example_config_freepdk45_row_addr_dff
* pin din_0
* pin dout_0
* pin din_1
* pin dout_1
* pin din_2
* pin dout_2
* pin din_3
* pin dout_3
* pin clk
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_row_addr_dff 1 2 3 4 5 6 7 8 9 10 11
* net 1 din_0
* net 2 dout_0
* net 3 din_1
* net 4 dout_1
* net 5 din_2
* net 6 dout_2
* net 7 din_3
* net 8 dout_3
* net 9 clk
* net 10 vdd
* net 11 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 9 10 11 dff
* cell instance $2 m0 *1 0,4.94
X$2 4 3 9 10 11 dff
* cell instance $3 r0 *1 0,4.94
X$3 6 5 9 10 11 dff
* cell instance $4 m0 *1 0,9.88
X$4 8 7 9 10 11 dff
.ENDS example_config_freepdk45_row_addr_dff

* cell example_config_freepdk45_control_logic_rw
* pin csb
* pin clk_buf
* pin clk
* pin web
* pin s_en
* pin w_en
* pin p_en_bar
* pin rbl_bl
* pin wl_en
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_control_logic_rw 1 2 4 8 13 15 16 17 18 19 20
* net 1 csb
* net 2 clk_buf
* net 4 clk
* net 8 web
* net 13 s_en
* net 15 w_en
* net 16 p_en_bar
* net 17 rbl_bl
* net 18 wl_en
* net 19 vdd
* net 20 gnd
* cell instance $1 r0 *1 0,0
X$1 1 3 8 10 5 2 19 20 example_config_freepdk45_dff_buf_array
* cell instance $3 m0 *1 6.385,4.94
X$3 2 6 19 20 example_config_freepdk45_pinv_3
* cell instance $4 r0 *1 6.385,4.94
X$4 9 2 3 19 20 example_config_freepdk45_pand2
* cell instance $11 r0 *1 6.385,0
X$11 2 4 19 20 example_config_freepdk45_pdriver_0
* cell instance $17 m0 *1 7.0725,4.94
X$17 7 6 3 19 20 example_config_freepdk45_pand2
* cell instance $20 r0 *1 6.385,9.88
X$20 15 5 12 7 19 20 example_config_freepdk45_pand3
* cell instance $24 m0 *1 6.385,9.88
X$24 13 11 7 10 19 20 example_config_freepdk45_pand3_0
* cell instance $25 m0 *1 6.385,19.76
X$25 18 7 19 20 example_config_freepdk45_pdriver_1
* cell instance $32 m0 *1 6.385,14.82
X$32 9 11 14 19 20 example_config_freepdk45_pnand2_1
* cell instance $40 m0 *1 0,32.11
X$40 11 17 19 20 example_config_freepdk45_delay_chain
* cell instance $41 r0 *1 6.385,14.82
X$41 11 12 19 20 example_config_freepdk45_pinv_3
* cell instance $52 m0 *1 7.2875,14.82
X$52 16 14 19 20 example_config_freepdk45_pdriver_4
.ENDS example_config_freepdk45_control_logic_rw

* cell example_config_freepdk45_bank
* pin din0_0
* pin din0_1
* pin w_en0
* pin p_en_bar0
* pin s_en0
* pin dout0_0
* pin dout0_1
* pin rbl_bl_0_0
* pin wl_en0
* pin addr0_0
* pin addr0_1
* pin addr0_2
* pin addr0_3
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_bank 1 2 3 4 5 6 7 8 14 20 21 22 23 36 37
* net 1 din0_0
* net 2 din0_1
* net 3 w_en0
* net 4 p_en_bar0
* net 5 s_en0
* net 6 dout0_0
* net 7 dout0_1
* net 8 rbl_bl_0_0
* net 14 wl_en0
* net 20 addr0_0
* net 21 addr0_1
* net 22 addr0_2
* net 23 addr0_3
* net 36 vdd
* net 37 gnd
* cell instance $1 m0 *1 10.49,13.04
X$1 4 5 3 10 11 12 13 1 2 6 7 8 9 36 37 example_config_freepdk45_port_data
* cell instance $5 r0 *1 10.49,13.04
X$5 15 17 16 18 19 25 27 24 8 9 10 11 12 13 30 26 28 31 33 29 34 32 35 36 37
+ example_config_freepdk45_capped_replica_bitcell_array
* cell instance $7 r0 *1 0,16.02
X$7 14 15 17 16 18 19 20 21 22 23 25 24 27 26 28 31 30 29 32 33 35 34 36 37
+ example_config_freepdk45_port_address
.ENDS example_config_freepdk45_bank

* cell example_config_freepdk45_pdriver_4
* pin Z
* pin A
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pdriver_4 1 2 4 5
* net 1 Z
* net 2 A
* net 4 vdd
* net 5 gnd
* cell instance $1 r0 *1 0.6875,0
X$1 3 1 4 5 example_config_freepdk45_pinv_5
* cell instance $2 r0 *1 0,0
X$2 2 3 4 5 example_config_freepdk45_pinv_5
.ENDS example_config_freepdk45_pdriver_4

* cell example_config_freepdk45_pnand2_1
* pin A
* pin B
* pin Z
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pnand2_1 1 2 3 4 5
* net 1 A
* net 2 B
* net 3 Z
* net 4 vdd
* net 5 gnd
* device instance $1 r0 *1 0.2325,2.21 PMOS_VTG
M$1 4 1 3 4 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.022275P PS=0.795U
+ PD=0.435U
* device instance $2 r0 *1 0.4475,2.21 PMOS_VTG
M$2 3 2 4 4 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.034425P PS=0.435U
+ PD=0.795U
* device instance $3 r0 *1 0.2325,0.215 NMOS_VTG
M$3 5 1 6 5 NMOS_VTG L=0.05U W=0.18U AS=0.02295P AD=0.01485P PS=0.615U PD=0.345U
* device instance $4 r0 *1 0.4475,0.215 NMOS_VTG
M$4 6 2 3 5 NMOS_VTG L=0.05U W=0.18U AS=0.01485P AD=0.02295P PS=0.345U PD=0.615U
.ENDS example_config_freepdk45_pnand2_1

* cell example_config_freepdk45_pand3_0
* pin Z
* pin A
* pin B
* pin C
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pand3_0 2 3 4 5 6 7
* net 2 Z
* net 3 A
* net 4 B
* net 5 C
* net 6 vdd
* net 7 gnd
* cell instance $1 r0 *1 0,0
X$1 3 4 5 1 6 7 example_config_freepdk45_pnand3_0
* cell instance $2 r0 *1 0.965,0
X$2 2 1 6 7 example_config_freepdk45_pdriver_3
.ENDS example_config_freepdk45_pand3_0

* cell example_config_freepdk45_pand3
* pin Z
* pin A
* pin B
* pin C
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pand3 2 3 4 5 6 7
* net 2 Z
* net 3 A
* net 4 B
* net 5 C
* net 6 vdd
* net 7 gnd
* cell instance $1 r0 *1 0.965,0
X$1 2 1 6 7 example_config_freepdk45_pdriver_2
* cell instance $2 r0 *1 0,0
X$2 3 4 5 1 6 7 example_config_freepdk45_pnand3_0
.ENDS example_config_freepdk45_pand3

* cell example_config_freepdk45_pdriver_0
* pin Z
* pin A
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pdriver_0 4 5 6 7
* net 4 Z
* net 5 A
* net 6 vdd
* net 7 gnd
* cell instance $1 r0 *1 0,0
X$1 5 1 6 7 example_config_freepdk45_pinv_5
* cell instance $2 r0 *1 0.6875,0
X$2 1 2 6 7 example_config_freepdk45_pinv_6
* cell instance $3 r0 *1 1.375,0
X$3 2 3 6 7 example_config_freepdk45_pinv_7
* cell instance $4 r0 *1 2.3375,0
X$4 3 4 6 7 example_config_freepdk45_pinv_8
.ENDS example_config_freepdk45_pdriver_0

* cell example_config_freepdk45_pand2
* pin Z
* pin A
* pin B
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pand2 2 3 4 5 6
* net 2 Z
* net 3 A
* net 4 B
* net 5 vdd
* net 6 gnd
* cell instance $1 r0 *1 0,0
X$1 3 4 1 5 6 example_config_freepdk45_pnand2_0
* cell instance $2 r0 *1 0.75,0
X$2 2 1 5 6 example_config_freepdk45_pdriver
.ENDS example_config_freepdk45_pand2

* cell example_config_freepdk45_dff_buf_array
* pin din_0
* pin dout_bar_0
* pin din_1
* pin dout_1
* pin dout_bar_1
* pin clk
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_dff_buf_array 1 3 4 5 6 7 8 9
* net 1 din_0
* net 2 dout_0
* net 3 dout_bar_0
* net 4 din_1
* net 5 dout_1
* net 6 dout_bar_1
* net 7 clk
* net 8 vdd
* net 9 gnd
* cell instance $1 r0 *1 0,0
X$1 3 2 7 1 8 9 example_config_freepdk45_dff_buf_0
* cell instance $2 m0 *1 0,4.94
X$2 6 5 7 4 8 9 example_config_freepdk45_dff_buf_0
.ENDS example_config_freepdk45_dff_buf_array

* cell example_config_freepdk45_pdriver_1
* pin Z
* pin A
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pdriver_1 2 3 4 5
* net 2 Z
* net 3 A
* net 4 vdd
* net 5 gnd
* cell instance $1 r0 *1 0.6875,0
X$1 1 2 4 5 example_config_freepdk45_pinv_7
* cell instance $2 r0 *1 0,0
X$2 3 1 4 5 example_config_freepdk45_pinv_5
.ENDS example_config_freepdk45_pdriver_1

* cell example_config_freepdk45_delay_chain
* pin out
* pin in
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_delay_chain 1 10 11 12
* net 1 out
* net 10 in
* net 11 vdd
* net 12 gnd
* cell instance $2 r0 *1 0.6875,19.76
X$2 1 37 11 12 example_config_freepdk45_pinv_10
* cell instance $5 r0 *1 1.375,19.76
X$5 1 36 11 12 example_config_freepdk45_pinv_10
* cell instance $8 r0 *1 2.0625,19.76
X$8 1 35 11 12 example_config_freepdk45_pinv_10
* cell instance $11 r0 *1 2.75,19.76
X$11 1 34 11 12 example_config_freepdk45_pinv_10
* cell instance $14 r0 *1 0,19.76
X$14 9 1 11 12 example_config_freepdk45_pinv_10
* cell instance $17 r0 *1 1.375,0
X$17 2 29 11 12 example_config_freepdk45_pinv_10
* cell instance $20 r0 *1 0.6875,0
X$20 2 46 11 12 example_config_freepdk45_pinv_10
* cell instance $23 m0 *1 0,4.94
X$23 2 3 11 12 example_config_freepdk45_pinv_10
* cell instance $25 r0 *1 2.0625,0
X$25 2 45 11 12 example_config_freepdk45_pinv_10
* cell instance $28 r0 *1 2.75,0
X$28 2 47 11 12 example_config_freepdk45_pinv_10
* cell instance $31 r0 *1 0,0
X$31 10 2 11 12 example_config_freepdk45_pinv_10
* cell instance $34 m0 *1 2.0625,4.94
X$34 3 22 11 12 example_config_freepdk45_pinv_10
* cell instance $37 r0 *1 0,4.94
X$37 3 4 11 12 example_config_freepdk45_pinv_10
* cell instance $39 m0 *1 2.75,4.94
X$39 3 23 11 12 example_config_freepdk45_pinv_10
* cell instance $42 m0 *1 0.6875,4.94
X$42 3 16 11 12 example_config_freepdk45_pinv_10
* cell instance $47 m0 *1 1.375,4.94
X$47 3 13 11 12 example_config_freepdk45_pinv_10
* cell instance $50 r0 *1 1.375,4.94
X$50 4 31 11 12 example_config_freepdk45_pinv_10
* cell instance $55 r0 *1 2.75,4.94
X$55 4 33 11 12 example_config_freepdk45_pinv_10
* cell instance $58 r0 *1 2.0625,4.94
X$58 4 32 11 12 example_config_freepdk45_pinv_10
* cell instance $61 m0 *1 0,9.88
X$61 4 5 11 12 example_config_freepdk45_pinv_10
* cell instance $63 r0 *1 0.6875,4.94
X$63 4 30 11 12 example_config_freepdk45_pinv_10
* cell instance $66 m0 *1 2.0625,9.88
X$66 5 15 11 12 example_config_freepdk45_pinv_10
* cell instance $69 r0 *1 0,9.88
X$69 5 6 11 12 example_config_freepdk45_pinv_10
* cell instance $71 m0 *1 0.6875,9.88
X$71 5 27 11 12 example_config_freepdk45_pinv_10
* cell instance $74 m0 *1 2.75,9.88
X$74 5 21 11 12 example_config_freepdk45_pinv_10
* cell instance $79 m0 *1 1.375,9.88
X$79 5 14 11 12 example_config_freepdk45_pinv_10
* cell instance $82 m0 *1 0,14.82
X$82 6 7 11 12 example_config_freepdk45_pinv_10
* cell instance $84 r0 *1 2.0625,9.88
X$84 6 43 11 12 example_config_freepdk45_pinv_10
* cell instance $87 r0 *1 0.6875,9.88
X$87 6 48 11 12 example_config_freepdk45_pinv_10
* cell instance $92 r0 *1 1.375,9.88
X$92 6 44 11 12 example_config_freepdk45_pinv_10
* cell instance $95 r0 *1 2.75,9.88
X$95 6 42 11 12 example_config_freepdk45_pinv_10
* cell instance $100 m0 *1 2.75,14.82
X$100 7 24 11 12 example_config_freepdk45_pinv_10
* cell instance $103 m0 *1 2.0625,14.82
X$103 7 25 11 12 example_config_freepdk45_pinv_10
* cell instance $106 m0 *1 0.6875,14.82
X$106 7 28 11 12 example_config_freepdk45_pinv_10
* cell instance $109 m0 *1 1.375,14.82
X$109 7 26 11 12 example_config_freepdk45_pinv_10
* cell instance $112 r0 *1 0,14.82
X$112 7 8 11 12 example_config_freepdk45_pinv_10
* cell instance $114 r0 *1 1.375,14.82
X$114 8 40 11 12 example_config_freepdk45_pinv_10
* cell instance $117 r0 *1 0.6875,14.82
X$117 8 41 11 12 example_config_freepdk45_pinv_10
* cell instance $120 r0 *1 2.0625,14.82
X$120 8 39 11 12 example_config_freepdk45_pinv_10
* cell instance $123 r0 *1 2.75,14.82
X$123 8 38 11 12 example_config_freepdk45_pinv_10
* cell instance $128 m0 *1 0,19.76
X$128 8 9 11 12 example_config_freepdk45_pinv_10
* cell instance $130 m0 *1 1.375,19.76
X$130 9 19 11 12 example_config_freepdk45_pinv_10
* cell instance $133 m0 *1 0.6875,19.76
X$133 9 20 11 12 example_config_freepdk45_pinv_10
* cell instance $136 m0 *1 2.0625,19.76
X$136 9 18 11 12 example_config_freepdk45_pinv_10
* cell instance $139 m0 *1 2.75,19.76
X$139 9 17 11 12 example_config_freepdk45_pinv_10
.ENDS example_config_freepdk45_delay_chain

* cell example_config_freepdk45_pinv_3
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pinv_3 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.17 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.09U AS=0.011475P AD=0.011475P PS=0.435U
+ PD=0.435U
* device instance $2 r0 *1 0.2325,2.21 PMOS_VTG
M$2 3 1 2 3 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.034425P PS=0.795U
+ PD=0.795U
.ENDS example_config_freepdk45_pinv_3

* cell example_config_freepdk45_port_address
* pin wl_en
* pin rbl_wl
* pin wl_0
* pin wl_1
* pin wl_2
* pin wl_3
* pin addr_0
* pin addr_1
* pin addr_2
* pin addr_3
* pin wl_4
* pin wl_5
* pin wl_6
* pin wl_7
* pin wl_8
* pin wl_9
* pin wl_10
* pin wl_11
* pin wl_13
* pin wl_12
* pin wl_15
* pin wl_14
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_port_address 1 2 5 7 9 10 11 12 13 14 16 18 21
+ 22 25 27 29 30 33 34 37 38 39 40
* net 1 wl_en
* net 2 rbl_wl
* net 5 wl_0
* net 7 wl_1
* net 9 wl_2
* net 10 wl_3
* net 11 addr_0
* net 12 addr_1
* net 13 addr_2
* net 14 addr_3
* net 16 wl_4
* net 18 wl_5
* net 21 wl_6
* net 22 wl_7
* net 25 wl_8
* net 27 wl_9
* net 29 wl_10
* net 30 wl_11
* net 33 wl_13
* net 34 wl_12
* net 37 wl_15
* net 38 wl_14
* net 39 vdd
* net 40 gnd
* cell instance $1 r0 *1 7.33,0
X$1 4 5 3 7 6 9 8 10 15 16 17 18 20 21 19 22 24 25 23 27 26 29 28 30 31 34 32
+ 33 35 38 36 37 1 39 40 example_config_freepdk45_wordline_driver_array
* cell instance $3 m0 *1 7.89,0
X$3 2 1 39 39 40 example_config_freepdk45_and2_dec_0
* cell instance $4 r0 *1 0,0
X$4 4 3 11 12 6 13 14 8 15 17 20 19 24 23 26 28 32 31 35 36 39 40
+ example_config_freepdk45_hierarchical_decoder
.ENDS example_config_freepdk45_port_address

* cell example_config_freepdk45_port_data
* pin p_en_bar
* pin s_en
* pin w_en
* pin bl_0
* pin br_0
* pin bl_1
* pin br_1
* pin din_0
* pin din_1
* pin dout_0
* pin dout_1
* pin rbl_bl
* pin rbl_br
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_port_data 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15
* net 1 p_en_bar
* net 2 s_en
* net 3 w_en
* net 4 bl_0
* net 5 br_0
* net 6 bl_1
* net 7 br_1
* net 8 din_0
* net 9 din_1
* net 10 dout_0
* net 11 dout_1
* net 12 rbl_bl
* net 13 rbl_br
* net 14 vdd
* net 15 gnd
* cell instance $1 m0 *1 0,1.845
X$1 1 12 13 4 5 6 7 14 example_config_freepdk45_precharge_array
* cell instance $2 m0 *1 0,8.36
X$2 2 4 5 10 6 7 11 14 15 example_config_freepdk45_sense_amp_array
* cell instance $3 m0 *1 0,13.04
X$3 3 8 4 5 9 6 7 14 15 example_config_freepdk45_write_driver_array
.ENDS example_config_freepdk45_port_data

* cell example_config_freepdk45_capped_replica_bitcell_array
* pin rbl_wl_0_0
* pin wl_0_0
* pin wl_0_1
* pin wl_0_2
* pin wl_0_3
* pin wl_0_4
* pin wl_0_6
* pin wl_0_5
* pin rbl_bl_0_0
* pin rbl_br_0_0
* pin bl_0_0
* pin br_0_0
* pin bl_0_1
* pin br_0_1
* pin wl_0_10
* pin wl_0_7
* pin wl_0_8
* pin wl_0_9
* pin wl_0_12
* pin wl_0_11
* pin wl_0_14
* pin wl_0_13
* pin wl_0_15
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_capped_replica_bitcell_array 1 2 3 4 5 6 7 8 9
+ 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25
* net 1 rbl_wl_0_0
* net 2 wl_0_0
* net 3 wl_0_1
* net 4 wl_0_2
* net 5 wl_0_3
* net 6 wl_0_4
* net 7 wl_0_6
* net 8 wl_0_5
* net 9 rbl_bl_0_0
* net 10 rbl_br_0_0
* net 11 bl_0_0
* net 12 br_0_0
* net 13 bl_0_1
* net 14 br_0_1
* net 15 wl_0_10
* net 16 wl_0_7
* net 17 wl_0_8
* net 18 wl_0_9
* net 19 wl_0_12
* net 20 wl_0_11
* net 21 wl_0_14
* net 22 wl_0_13
* net 23 wl_0_15
* net 24 vdd
* net 25 gnd
* cell instance $1 r0 *1 1.64,1.615
X$1 1 9 10 11 12 13 14 2 3 4 5 6 8 7 16 17 18 15 20 19 22 21 23 24 25
+ example_config_freepdk45_replica_bitcell_array
* cell instance $2 r0 *1 0.935,0.25
X$2 25 1 2 3 4 5 6 8 7 16 17 18 15 20 19 22 21 23 25 24 25
+ example_config_freepdk45_dummy_array_2
* cell instance $3 r0 *1 3.755,0.25
X$3 25 1 2 3 4 5 6 8 7 16 17 18 15 20 19 22 21 23 25 24 25
+ example_config_freepdk45_dummy_array_3
* cell instance $4 r0 *1 1.64,0.25
X$4 25 24 25 example_config_freepdk45_dummy_array_1
* cell instance $5 r0 *1 1.64,24.82
X$5 25 24 25 example_config_freepdk45_dummy_array_0
.ENDS example_config_freepdk45_capped_replica_bitcell_array

* cell example_config_freepdk45_pdriver_3
* pin Z
* pin A
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pdriver_3 1 2 3 4
* net 1 Z
* net 2 A
* net 3 vdd
* net 4 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 3 4 example_config_freepdk45_pinv_6
.ENDS example_config_freepdk45_pdriver_3

* cell example_config_freepdk45_pdriver_2
* pin Z
* pin A
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pdriver_2 1 2 3 4
* net 1 Z
* net 2 A
* net 3 vdd
* net 4 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 3 4 example_config_freepdk45_pinv_9
.ENDS example_config_freepdk45_pdriver_2

* cell example_config_freepdk45_pnand3_0
* pin A
* pin B
* pin C
* pin Z
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pnand3_0 1 2 3 4 5 6
* net 1 A
* net 2 B
* net 3 C
* net 4 Z
* net 5 vdd
* net 6 gnd
* device instance $1 r0 *1 0.2325,2.21 PMOS_VTG
M$1 5 1 4 5 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.022275P PS=0.795U
+ PD=0.435U
* device instance $2 r0 *1 0.4475,2.21 PMOS_VTG
M$2 4 2 5 5 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.022275P PS=0.435U
+ PD=0.435U
* device instance $3 r0 *1 0.6625,2.21 PMOS_VTG
M$3 5 3 4 5 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.034425P PS=0.435U
+ PD=0.795U
* device instance $4 r0 *1 0.2325,0.215 NMOS_VTG
M$4 6 1 8 6 NMOS_VTG L=0.05U W=0.18U AS=0.02295P AD=0.01485P PS=0.615U PD=0.345U
* device instance $5 r0 *1 0.4475,0.215 NMOS_VTG
M$5 8 2 7 6 NMOS_VTG L=0.05U W=0.18U AS=0.01485P AD=0.01485P PS=0.345U PD=0.345U
* device instance $6 r0 *1 0.6625,0.215 NMOS_VTG
M$6 7 3 4 6 NMOS_VTG L=0.05U W=0.18U AS=0.01485P AD=0.02295P PS=0.345U PD=0.615U
.ENDS example_config_freepdk45_pnand3_0

* cell example_config_freepdk45_pinv_8
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pinv_8 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.26 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=1.35U AS=0.155925P AD=0.155925P PS=2.775U
+ PD=2.775U
* device instance $6 r0 *1 0.2325,1.94 PMOS_VTG
M$6 3 1 2 3 PMOS_VTG L=0.05U W=4.05U AS=0.467775P AD=0.467775P PS=6.015U
+ PD=6.015U
.ENDS example_config_freepdk45_pinv_8

* cell example_config_freepdk45_pdriver
* pin Z
* pin A
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pdriver 1 2 3 4
* net 1 Z
* net 2 A
* net 3 vdd
* net 4 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 3 4 example_config_freepdk45_pinv_2
.ENDS example_config_freepdk45_pdriver

* cell example_config_freepdk45_pnand2_0
* pin A
* pin B
* pin Z
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pnand2_0 1 2 3 4 5
* net 1 A
* net 2 B
* net 3 Z
* net 4 vdd
* net 5 gnd
* device instance $1 r0 *1 0.2325,2.21 PMOS_VTG
M$1 4 1 3 4 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.022275P PS=0.795U
+ PD=0.435U
* device instance $2 r0 *1 0.4475,2.21 PMOS_VTG
M$2 3 2 4 4 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.034425P PS=0.435U
+ PD=0.795U
* device instance $3 r0 *1 0.2325,0.215 NMOS_VTG
M$3 5 1 6 5 NMOS_VTG L=0.05U W=0.18U AS=0.02295P AD=0.01485P PS=0.615U PD=0.345U
* device instance $4 r0 *1 0.4475,0.215 NMOS_VTG
M$4 6 2 3 5 NMOS_VTG L=0.05U W=0.18U AS=0.01485P AD=0.02295P PS=0.345U PD=0.615U
.ENDS example_config_freepdk45_pnand2_0

* cell example_config_freepdk45_dff_buf_0
* pin Qb
* pin Q
* pin clk
* pin D
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_dff_buf_0 1 2 4 5 6 7
* net 1 Qb
* net 2 Q
* net 4 clk
* net 5 D
* net 6 vdd
* net 7 gnd
* cell instance $1 r0 *1 3.195,0
X$1 3 1 6 7 example_config_freepdk45_pinv_0
* cell instance $2 r0 *1 3.8825,0
X$2 1 2 6 7 example_config_freepdk45_pinv_1
* cell instance $5 r0 *1 0,0
X$5 3 5 4 6 7 dff
.ENDS example_config_freepdk45_dff_buf_0

* cell example_config_freepdk45_pinv_7
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pinv_7 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.2375 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.45U AS=0.054P AD=0.054P PS=1.155U PD=1.155U
* device instance $3 r0 *1 0.2325,2.0075 PMOS_VTG
M$3 3 1 2 3 PMOS_VTG L=0.05U W=1.35U AS=0.162P AD=0.162P PS=2.505U PD=2.505U
.ENDS example_config_freepdk45_pinv_7

* cell example_config_freepdk45_pinv_5
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pinv_5 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.17 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.09U AS=0.011475P AD=0.011475P PS=0.435U
+ PD=0.435U
* device instance $2 r0 *1 0.2325,2.21 PMOS_VTG
M$2 3 1 2 3 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.034425P PS=0.795U
+ PD=0.795U
.ENDS example_config_freepdk45_pinv_5

* cell example_config_freepdk45_pinv_10
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pinv_10 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.17 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.09U AS=0.011475P AD=0.011475P PS=0.435U
+ PD=0.435U
* device instance $2 r0 *1 0.2325,2.21 PMOS_VTG
M$2 3 1 2 3 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.034425P PS=0.795U
+ PD=0.795U
.ENDS example_config_freepdk45_pinv_10

* cell example_config_freepdk45_and2_dec_0
* pin Z
* pin A
* pin B
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_and2_dec_0 2 3 4 5 6
* net 2 Z
* net 3 A
* net 4 B
* net 5 vdd
* net 6 gnd
* cell instance $1 r0 *1 0.9025,0
X$1 1 2 5 6 example_config_freepdk45_pinv
* cell instance $2 r0 *1 0,0
X$2 3 4 1 5 6 example_config_freepdk45_pnand2
.ENDS example_config_freepdk45_and2_dec_0

* cell example_config_freepdk45_wordline_driver_array
* pin in_0
* pin wl_0
* pin in_1
* pin wl_1
* pin in_2
* pin wl_2
* pin in_3
* pin wl_3
* pin in_4
* pin wl_4
* pin in_5
* pin wl_5
* pin in_6
* pin wl_6
* pin in_7
* pin wl_7
* pin in_8
* pin wl_8
* pin in_9
* pin wl_9
* pin in_10
* pin wl_10
* pin in_11
* pin wl_11
* pin in_12
* pin wl_12
* pin in_13
* pin wl_13
* pin in_14
* pin wl_14
* pin in_15
* pin wl_15
* pin en
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_wordline_driver_array 1 2 3 4 5 6 7 8 9 10 11
+ 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35
* net 1 in_0
* net 2 wl_0
* net 3 in_1
* net 4 wl_1
* net 5 in_2
* net 6 wl_2
* net 7 in_3
* net 8 wl_3
* net 9 in_4
* net 10 wl_4
* net 11 in_5
* net 12 wl_5
* net 13 in_6
* net 14 wl_6
* net 15 in_7
* net 16 wl_7
* net 17 in_8
* net 18 wl_8
* net 19 in_9
* net 20 wl_9
* net 21 in_10
* net 22 wl_10
* net 23 in_11
* net 24 wl_11
* net 25 in_12
* net 26 wl_12
* net 27 in_13
* net 28 wl_13
* net 29 in_14
* net 30 wl_14
* net 31 in_15
* net 32 wl_15
* net 33 en
* net 34 vdd
* net 35 gnd
* cell instance $1 r0 *1 0.56,0
X$1 2 1 33 34 35 example_config_freepdk45_wordline_driver
* cell instance $2 m0 *1 0.56,2.73
X$2 4 3 33 34 35 example_config_freepdk45_wordline_driver
* cell instance $3 r0 *1 0.56,2.73
X$3 6 5 33 34 35 example_config_freepdk45_wordline_driver
* cell instance $4 m0 *1 0.56,5.46
X$4 8 7 33 34 35 example_config_freepdk45_wordline_driver
* cell instance $5 r0 *1 0.56,5.46
X$5 10 9 33 34 35 example_config_freepdk45_wordline_driver
* cell instance $6 m0 *1 0.56,8.19
X$6 12 11 33 34 35 example_config_freepdk45_wordline_driver
* cell instance $7 r0 *1 0.56,8.19
X$7 14 13 33 34 35 example_config_freepdk45_wordline_driver
* cell instance $8 m0 *1 0.56,10.92
X$8 16 15 33 34 35 example_config_freepdk45_wordline_driver
* cell instance $9 r0 *1 0.56,10.92
X$9 18 17 33 34 35 example_config_freepdk45_wordline_driver
* cell instance $10 m0 *1 0.56,13.65
X$10 20 19 33 34 35 example_config_freepdk45_wordline_driver
* cell instance $11 r0 *1 0.56,13.65
X$11 22 21 33 34 35 example_config_freepdk45_wordline_driver
* cell instance $12 m0 *1 0.56,16.38
X$12 24 23 33 34 35 example_config_freepdk45_wordline_driver
* cell instance $13 r0 *1 0.56,16.38
X$13 26 25 33 34 35 example_config_freepdk45_wordline_driver
* cell instance $14 m0 *1 0.56,19.11
X$14 28 27 33 34 35 example_config_freepdk45_wordline_driver
* cell instance $15 r0 *1 0.56,19.11
X$15 30 29 33 34 35 example_config_freepdk45_wordline_driver
* cell instance $16 m0 *1 0.56,21.84
X$16 32 31 33 34 35 example_config_freepdk45_wordline_driver
.ENDS example_config_freepdk45_wordline_driver_array

* cell example_config_freepdk45_hierarchical_decoder
* pin decode_0
* pin decode_1
* pin addr_0
* pin addr_1
* pin decode_2
* pin addr_2
* pin addr_3
* pin decode_3
* pin decode_4
* pin decode_5
* pin decode_6
* pin decode_7
* pin decode_8
* pin decode_9
* pin decode_10
* pin decode_11
* pin decode_13
* pin decode_12
* pin decode_14
* pin decode_15
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_hierarchical_decoder 4 5 6 7 10 11 12 14 15 16
+ 17 19 21 22 23 24 25 26 27 28 29 30
* net 4 decode_0
* net 5 decode_1
* net 6 addr_0
* net 7 addr_1
* net 10 decode_2
* net 11 addr_2
* net 12 addr_3
* net 14 decode_3
* net 15 decode_4
* net 16 decode_5
* net 17 decode_6
* net 19 decode_7
* net 21 decode_8
* net 22 decode_9
* net 23 decode_10
* net 24 decode_11
* net 25 decode_13
* net 26 decode_12
* net 27 decode_14
* net 28 decode_15
* net 29 vdd
* net 30 gnd
* cell instance $2 r0 *1 5.74,10.92
X$2 21 1 18 29 30 example_config_freepdk45_and2_dec
* cell instance $3 r0 *1 5.74,5.46
X$3 15 1 13 29 30 example_config_freepdk45_and2_dec
* cell instance $4 r0 *1 5.74,0
X$4 4 1 3 29 30 example_config_freepdk45_and2_dec
* cell instance $5 r0 *1 5.74,16.38
X$5 26 1 20 29 30 example_config_freepdk45_and2_dec
* cell instance $7 r0 *1 0.6625,0
X$7 6 7 1 2 9 8 29 30 example_config_freepdk45_hierarchical_predecode2x4
* cell instance $14 m0 *1 5.74,13.65
X$14 22 2 18 29 30 example_config_freepdk45_and2_dec
* cell instance $15 m0 *1 5.74,8.19
X$15 16 2 13 29 30 example_config_freepdk45_and2_dec
* cell instance $16 m0 *1 5.74,2.73
X$16 5 2 3 29 30 example_config_freepdk45_and2_dec
* cell instance $17 m0 *1 5.74,19.11
X$17 25 2 20 29 30 example_config_freepdk45_and2_dec
* cell instance $25 m0 *1 5.74,5.46
X$25 14 8 3 29 30 example_config_freepdk45_and2_dec
* cell instance $26 r0 *1 5.74,2.73
X$26 10 9 3 29 30 example_config_freepdk45_and2_dec
* cell instance $28 r0 *1 0.6625,8.19
X$28 11 12 3 13 18 20 29 30 example_config_freepdk45_hierarchical_predecode2x4
* cell instance $39 m0 *1 5.74,16.38
X$39 24 8 18 29 30 example_config_freepdk45_and2_dec
* cell instance $40 m0 *1 5.74,21.84
X$40 28 8 20 29 30 example_config_freepdk45_and2_dec
* cell instance $41 m0 *1 5.74,10.92
X$41 19 8 13 29 30 example_config_freepdk45_and2_dec
* cell instance $49 r0 *1 5.74,8.19
X$49 17 9 13 29 30 example_config_freepdk45_and2_dec
* cell instance $50 r0 *1 5.74,13.65
X$50 23 9 18 29 30 example_config_freepdk45_and2_dec
* cell instance $51 r0 *1 5.74,19.11
X$51 27 9 20 29 30 example_config_freepdk45_and2_dec
.ENDS example_config_freepdk45_hierarchical_decoder

* cell example_config_freepdk45_write_driver_array
* pin en
* pin data_0
* pin bl_0
* pin br_0
* pin data_1
* pin bl_1
* pin br_1
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_write_driver_array 1 2 3 4 5 6 7 8 9
* net 1 en
* net 2 data_0
* net 3 bl_0
* net 4 br_0
* net 5 data_1
* net 6 bl_1
* net 7 br_1
* net 8 vdd
* net 9 gnd
* cell instance $1 r0 *1 2.345,0
X$1 2 1 4 3 8 9 write_driver
* cell instance $2 r0 *1 3.05,0
X$2 5 1 7 6 8 9 write_driver
.ENDS example_config_freepdk45_write_driver_array

* cell example_config_freepdk45_sense_amp_array
* pin en
* pin bl_0
* pin br_0
* pin data_0
* pin bl_1
* pin br_1
* pin data_1
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_sense_amp_array 1 2 3 4 5 6 7 8 9
* net 1 en
* net 2 bl_0
* net 3 br_0
* net 4 data_0
* net 5 bl_1
* net 6 br_1
* net 7 data_1
* net 8 vdd
* net 9 gnd
* cell instance $1 r0 *1 3.05,0
X$1 6 7 5 1 8 9 sense_amp
* cell instance $2 r0 *1 2.345,0
X$2 3 4 2 1 8 9 sense_amp
.ENDS example_config_freepdk45_sense_amp_array

* cell example_config_freepdk45_precharge_array
* pin en_bar
* pin bl_0
* pin br_0
* pin bl_1
* pin br_1
* pin bl_2
* pin br_2
* pin vdd
.SUBCKT example_config_freepdk45_precharge_array 1 2 3 4 5 6 7 8
* net 1 en_bar
* net 2 bl_0
* net 3 br_0
* net 4 bl_1
* net 5 br_1
* net 6 bl_2
* net 7 br_2
* net 8 vdd
* cell instance $1 r0 *1 2.345,0
X$1 1 4 5 8 example_config_freepdk45_precharge_0
* cell instance $2 r0 *1 1.64,0
X$2 1 2 3 8 example_config_freepdk45_precharge_0
* cell instance $3 r0 *1 3.05,0
X$3 1 6 7 8 example_config_freepdk45_precharge_0
.ENDS example_config_freepdk45_precharge_array

* cell example_config_freepdk45_dummy_array_1
* pin wl_0_0
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_dummy_array_1 1 2 3
* net 1 wl_0_0
* net 2 vdd
* net 3 gnd
* cell instance $1 r0 *1 0,0
X$1 1 2 3 dummy_cell_1rw
* cell instance $2 r0 *1 0.705,0
X$2 1 2 3 dummy_cell_1rw
* cell instance $3 r0 *1 1.41,0
X$3 1 2 3 dummy_cell_1rw
.ENDS example_config_freepdk45_dummy_array_1

* cell example_config_freepdk45_dummy_array_0
* pin wl_0_0
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_dummy_array_0 1 2 3
* net 1 wl_0_0
* net 2 vdd
* net 3 gnd
* cell instance $1 r0 *1 0,0
X$1 1 2 3 dummy_cell_1rw
* cell instance $2 r0 *1 0.705,0
X$2 1 2 3 dummy_cell_1rw
* cell instance $3 r0 *1 1.41,0
X$3 1 2 3 dummy_cell_1rw
.ENDS example_config_freepdk45_dummy_array_0

* cell example_config_freepdk45_dummy_array_3
* pin wl_0_0
* pin wl_0_1
* pin wl_0_2
* pin wl_0_3
* pin wl_0_4
* pin wl_0_5
* pin wl_0_6
* pin wl_0_7
* pin wl_0_8
* pin wl_0_9
* pin wl_0_10
* pin wl_0_11
* pin wl_0_12
* pin wl_0_13
* pin wl_0_14
* pin wl_0_15
* pin wl_0_16
* pin wl_0_17
* pin wl_0_18
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_dummy_array_3 1 2 3 4 5 6 7 8 9 10 11 12 13 14
+ 15 16 17 18 19 20 21
* net 1 wl_0_0
* net 2 wl_0_1
* net 3 wl_0_2
* net 4 wl_0_3
* net 5 wl_0_4
* net 6 wl_0_5
* net 7 wl_0_6
* net 8 wl_0_7
* net 9 wl_0_8
* net 10 wl_0_9
* net 11 wl_0_10
* net 12 wl_0_11
* net 13 wl_0_12
* net 14 wl_0_13
* net 15 wl_0_14
* net 16 wl_0_15
* net 17 wl_0_16
* net 18 wl_0_17
* net 19 wl_0_18
* net 20 vdd
* net 21 gnd
* cell instance $1 r0 *1 0,0
X$1 1 20 21 dummy_cell_1rw
* cell instance $2 m0 *1 0,2.73
X$2 2 20 21 dummy_cell_1rw
* cell instance $3 r0 *1 0,2.73
X$3 3 20 21 dummy_cell_1rw
* cell instance $4 m0 *1 0,5.46
X$4 4 20 21 dummy_cell_1rw
* cell instance $5 r0 *1 0,5.46
X$5 5 20 21 dummy_cell_1rw
* cell instance $6 m0 *1 0,8.19
X$6 6 20 21 dummy_cell_1rw
* cell instance $7 r0 *1 0,8.19
X$7 7 20 21 dummy_cell_1rw
* cell instance $8 m0 *1 0,10.92
X$8 8 20 21 dummy_cell_1rw
* cell instance $9 r0 *1 0,10.92
X$9 9 20 21 dummy_cell_1rw
* cell instance $10 m0 *1 0,13.65
X$10 10 20 21 dummy_cell_1rw
* cell instance $11 r0 *1 0,13.65
X$11 11 20 21 dummy_cell_1rw
* cell instance $12 m0 *1 0,16.38
X$12 12 20 21 dummy_cell_1rw
* cell instance $13 r0 *1 0,16.38
X$13 13 20 21 dummy_cell_1rw
* cell instance $14 m0 *1 0,19.11
X$14 14 20 21 dummy_cell_1rw
* cell instance $15 r0 *1 0,19.11
X$15 15 20 21 dummy_cell_1rw
* cell instance $16 m0 *1 0,21.84
X$16 16 20 21 dummy_cell_1rw
* cell instance $17 r0 *1 0,21.84
X$17 17 20 21 dummy_cell_1rw
* cell instance $18 m0 *1 0,24.57
X$18 18 20 21 dummy_cell_1rw
* cell instance $19 r0 *1 0,24.57
X$19 19 20 21 dummy_cell_1rw
.ENDS example_config_freepdk45_dummy_array_3

* cell example_config_freepdk45_dummy_array_2
* pin wl_0_0
* pin wl_0_1
* pin wl_0_2
* pin wl_0_3
* pin wl_0_4
* pin wl_0_5
* pin wl_0_6
* pin wl_0_7
* pin wl_0_8
* pin wl_0_9
* pin wl_0_10
* pin wl_0_11
* pin wl_0_12
* pin wl_0_13
* pin wl_0_14
* pin wl_0_15
* pin wl_0_16
* pin wl_0_17
* pin wl_0_18
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_dummy_array_2 1 2 3 4 5 6 7 8 9 10 11 12 13 14
+ 15 16 17 18 19 20 21
* net 1 wl_0_0
* net 2 wl_0_1
* net 3 wl_0_2
* net 4 wl_0_3
* net 5 wl_0_4
* net 6 wl_0_5
* net 7 wl_0_6
* net 8 wl_0_7
* net 9 wl_0_8
* net 10 wl_0_9
* net 11 wl_0_10
* net 12 wl_0_11
* net 13 wl_0_12
* net 14 wl_0_13
* net 15 wl_0_14
* net 16 wl_0_15
* net 17 wl_0_16
* net 18 wl_0_17
* net 19 wl_0_18
* net 20 vdd
* net 21 gnd
* cell instance $1 r0 *1 0,0
X$1 1 20 21 dummy_cell_1rw
* cell instance $2 m0 *1 0,2.73
X$2 2 20 21 dummy_cell_1rw
* cell instance $3 r0 *1 0,2.73
X$3 3 20 21 dummy_cell_1rw
* cell instance $4 m0 *1 0,5.46
X$4 4 20 21 dummy_cell_1rw
* cell instance $5 r0 *1 0,5.46
X$5 5 20 21 dummy_cell_1rw
* cell instance $6 m0 *1 0,8.19
X$6 6 20 21 dummy_cell_1rw
* cell instance $7 r0 *1 0,8.19
X$7 7 20 21 dummy_cell_1rw
* cell instance $8 m0 *1 0,10.92
X$8 8 20 21 dummy_cell_1rw
* cell instance $9 r0 *1 0,10.92
X$9 9 20 21 dummy_cell_1rw
* cell instance $10 m0 *1 0,13.65
X$10 10 20 21 dummy_cell_1rw
* cell instance $11 r0 *1 0,13.65
X$11 11 20 21 dummy_cell_1rw
* cell instance $12 m0 *1 0,16.38
X$12 12 20 21 dummy_cell_1rw
* cell instance $13 r0 *1 0,16.38
X$13 13 20 21 dummy_cell_1rw
* cell instance $14 m0 *1 0,19.11
X$14 14 20 21 dummy_cell_1rw
* cell instance $15 r0 *1 0,19.11
X$15 15 20 21 dummy_cell_1rw
* cell instance $16 m0 *1 0,21.84
X$16 16 20 21 dummy_cell_1rw
* cell instance $17 r0 *1 0,21.84
X$17 17 20 21 dummy_cell_1rw
* cell instance $18 m0 *1 0,24.57
X$18 18 20 21 dummy_cell_1rw
* cell instance $19 r0 *1 0,24.57
X$19 19 20 21 dummy_cell_1rw
.ENDS example_config_freepdk45_dummy_array_2

* cell example_config_freepdk45_replica_bitcell_array
* pin rbl_wl_0_0
* pin rbl_bl_0_0
* pin rbl_br_0_0
* pin bl_0_0
* pin br_0_0
* pin bl_0_1
* pin br_0_1
* pin wl_0_0
* pin wl_0_1
* pin wl_0_2
* pin wl_0_3
* pin wl_0_4
* pin wl_0_5
* pin wl_0_6
* pin wl_0_7
* pin wl_0_8
* pin wl_0_9
* pin wl_0_10
* pin wl_0_11
* pin wl_0_12
* pin wl_0_13
* pin wl_0_14
* pin wl_0_15
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_replica_bitcell_array 1 2 3 4 5 6 7 8 9 10 11
+ 12 13 14 15 16 17 18 19 20 21 22 23 24 25
* net 1 rbl_wl_0_0
* net 2 rbl_bl_0_0
* net 3 rbl_br_0_0
* net 4 bl_0_0
* net 5 br_0_0
* net 6 bl_0_1
* net 7 br_0_1
* net 8 wl_0_0
* net 9 wl_0_1
* net 10 wl_0_2
* net 11 wl_0_3
* net 12 wl_0_4
* net 13 wl_0_5
* net 14 wl_0_6
* net 15 wl_0_7
* net 16 wl_0_8
* net 17 wl_0_9
* net 18 wl_0_10
* net 19 wl_0_11
* net 20 wl_0_12
* net 21 wl_0_13
* net 22 wl_0_14
* net 23 wl_0_15
* net 24 vdd
* net 25 gnd
* cell instance $1 r0 *1 0,0
X$1 1 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 2 3 24 25
+ example_config_freepdk45_replica_column
* cell instance $2 m0 *1 0.705,1.365
X$2 1 24 25 example_config_freepdk45_dummy_array
* cell instance $3 r0 *1 0.705,1.365
X$3 8 9 10 11 12 13 14 15 4 5 6 7 16 17 18 19 20 21 22 23 24 25
+ example_config_freepdk45_bitcell_array
.ENDS example_config_freepdk45_replica_bitcell_array

* cell example_config_freepdk45_pinv_9
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pinv_9 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.275 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.9U AS=0.10575P AD=0.10575P PS=1.905U PD=1.905U
* device instance $4 r0 *1 0.2325,1.895 PMOS_VTG
M$4 3 1 2 3 PMOS_VTG L=0.05U W=2.7U AS=0.31725P AD=0.31725P PS=4.305U PD=4.305U
.ENDS example_config_freepdk45_pinv_9

* cell example_config_freepdk45_pinv_6
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pinv_6 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.215 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.18U AS=0.02295P AD=0.02295P PS=0.615U PD=0.615U
* device instance $2 r0 *1 0.2325,2.075 PMOS_VTG
M$2 3 1 2 3 PMOS_VTG L=0.05U W=0.54U AS=0.06885P AD=0.06885P PS=1.335U PD=1.335U
.ENDS example_config_freepdk45_pinv_6

* cell example_config_freepdk45_pinv_2
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pinv_2 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.26 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=1.08U AS=0.12555P AD=0.12555P PS=2.28U PD=2.28U
* device instance $5 r0 *1 0.2325,1.94 PMOS_VTG
M$5 3 1 2 3 PMOS_VTG L=0.05U W=3.24U AS=0.37665P AD=0.37665P PS=4.98U PD=4.98U
.ENDS example_config_freepdk45_pinv_2

* cell example_config_freepdk45_pinv_1
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pinv_1 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.215 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.36U AS=0.0432P AD=0.0432P PS=1.02U PD=1.02U
* device instance $3 r0 *1 0.2325,2.075 PMOS_VTG
M$3 3 1 2 3 PMOS_VTG L=0.05U W=1.08U AS=0.1296P AD=0.1296P PS=2.1U PD=2.1U
.ENDS example_config_freepdk45_pinv_1

* cell example_config_freepdk45_pinv_0
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pinv_0 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.215 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.18U AS=0.02295P AD=0.02295P PS=0.615U PD=0.615U
* device instance $2 r0 *1 0.2325,2.075 PMOS_VTG
M$2 3 1 2 3 PMOS_VTG L=0.05U W=0.54U AS=0.06885P AD=0.06885P PS=1.335U PD=1.335U
.ENDS example_config_freepdk45_pinv_0

* cell dff
* pin Q
* pin D
* pin clk
* pin vdd
* pin gnd
.SUBCKT dff 2 5 7 16 17
* net 2 Q
* net 5 D
* net 7 clk
* net 16 vdd
* net 17 gnd
* device instance $1 r0 *1 0.2925,1.5425 PMOS_VTG
M$1 16 5 13 16 PMOS_VTG L=0.05U W=0.5U AS=0.0525P AD=0.035P PS=1.21U PD=0.64U
* device instance $2 r0 *1 0.4825,1.5425 PMOS_VTG
M$2 13 7 4 16 PMOS_VTG L=0.05U W=0.5U AS=0.035P AD=0.035P PS=0.64U PD=0.64U
* device instance $3 r0 *1 0.6725,1.5425 PMOS_VTG
M$3 4 1 14 16 PMOS_VTG L=0.05U W=0.5U AS=0.035P AD=0.035P PS=0.64U PD=0.64U
* device instance $4 r0 *1 0.8625,1.5425 PMOS_VTG
M$4 14 6 16 16 PMOS_VTG L=0.05U W=0.5U AS=0.035P AD=0.0851P PS=0.64U PD=1.275U
* device instance $5 r0 *1 1.1575,1.5425 PMOS_VTG
M$5 16 4 6 16 PMOS_VTG L=0.05U W=0.5U AS=0.0851P AD=0.0525P PS=1.275U PD=1.21U
* device instance $6 r0 *1 2.2325,1.4525 PMOS_VTG
M$6 8 7 12 16 PMOS_VTG L=0.05U W=0.25U AS=0.038125P AD=0.0375P PS=0.7U PD=0.8U
* device instance $7 r0 *1 1.7925,1.5775 PMOS_VTG
M$7 16 6 15 16 PMOS_VTG L=0.05U W=0.5U AS=0.0875P AD=0.035P PS=1.245U PD=0.64U
* device instance $8 r0 *1 1.9825,1.5775 PMOS_VTG
M$8 15 1 8 16 PMOS_VTG L=0.05U W=0.5U AS=0.035P AD=0.038125P PS=0.64U PD=0.7U
* device instance $9 r0 *1 1.4975,1.65 PMOS_VTG
M$9 1 7 16 16 PMOS_VTG L=0.05U W=1U AS=0.105P AD=0.0875P PS=2.21U PD=1.245U
* device instance $10 r0 *1 2.3225,2.0175 PMOS_VTG
M$10 16 2 12 16 PMOS_VTG L=0.05U W=0.25U AS=0.055125P AD=0.02625P PS=1.21U
+ PD=0.71U
* device instance $11 r0 *1 2.5825,1.7925 PMOS_VTG
M$11 16 8 2 16 PMOS_VTG L=0.05U W=1U AS=0.055125P AD=0.105P PS=1.21U PD=2.21U
* device instance $12 r0 *1 2.0475,0.3475 NMOS_VTG
M$12 17 2 3 17 NMOS_VTG L=0.05U W=0.25U AS=0.02625P AD=0.02625P PS=0.71U
+ PD=0.71U
* device instance $13 r0 *1 2.5825,0.7125 NMOS_VTG
M$13 17 8 2 17 NMOS_VTG L=0.05U W=0.5U AS=0.0775P AD=0.0525P PS=1.31U PD=1.21U
* device instance $14 r0 *1 0.2925,0.725 NMOS_VTG
M$14 17 5 9 17 NMOS_VTG L=0.05U W=0.25U AS=0.02625P AD=0.0175P PS=0.71U PD=0.39U
* device instance $15 r0 *1 0.4825,0.725 NMOS_VTG
M$15 9 1 4 17 NMOS_VTG L=0.05U W=0.25U AS=0.0175P AD=0.0175P PS=0.39U PD=0.39U
* device instance $16 r0 *1 0.6725,0.725 NMOS_VTG
M$16 4 7 10 17 NMOS_VTG L=0.05U W=0.25U AS=0.0175P AD=0.0175P PS=0.39U PD=0.39U
* device instance $17 r0 *1 0.8625,0.725 NMOS_VTG
M$17 17 6 10 17 NMOS_VTG L=0.05U W=0.25U AS=0.0502P AD=0.0175P PS=0.93U PD=0.39U
* device instance $18 r0 *1 1.1575,0.725 NMOS_VTG
M$18 17 4 6 17 NMOS_VTG L=0.05U W=0.25U AS=0.0502P AD=0.02625P PS=0.93U PD=0.71U
* device instance $19 r0 *1 1.4975,0.6575 NMOS_VTG
M$19 1 7 17 17 NMOS_VTG L=0.05U W=0.5U AS=0.0525P AD=0.04375P PS=1.21U PD=0.745U
* device instance $20 r0 *1 1.7925,0.7825 NMOS_VTG
M$20 17 6 11 17 NMOS_VTG L=0.05U W=0.25U AS=0.04375P AD=0.0175P PS=0.745U
+ PD=0.39U
* device instance $21 r0 *1 1.9825,0.7825 NMOS_VTG
M$21 11 7 8 17 NMOS_VTG L=0.05U W=0.25U AS=0.0175P AD=0.0175P PS=0.39U PD=0.39U
* device instance $22 r0 *1 2.1725,0.7825 NMOS_VTG
M$22 8 1 3 17 NMOS_VTG L=0.05U W=0.25U AS=0.0175P AD=0.0275P PS=0.39U PD=0.72U
.ENDS dff

* cell example_config_freepdk45_wordline_driver
* pin Z
* pin A
* pin B
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_wordline_driver 2 3 4 5 6
* net 2 Z
* net 3 A
* net 4 B
* net 5 vdd
* net 6 gnd
* cell instance $1 r0 *1 0.9025,0
X$1 1 2 5 6 example_config_freepdk45_pinv
* cell instance $2 r0 *1 0,0
X$2 3 4 1 5 6 example_config_freepdk45_pnand2
.ENDS example_config_freepdk45_wordline_driver

* cell example_config_freepdk45_hierarchical_predecode2x4
* pin in_0
* pin in_1
* pin out_0
* pin out_1
* pin out_2
* pin out_3
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_hierarchical_predecode2x4 1 2 5 6 7 8 9 10
* net 1 in_0
* net 2 in_1
* net 5 out_0
* net 6 out_1
* net 7 out_2
* net 8 out_3
* net 9 vdd
* net 10 gnd
* cell instance $1 m0 *1 2.0875,5.46
X$1 8 1 2 9 10 example_config_freepdk45_and2_dec
* cell instance $2 m0 *1 2.0875,2.73
X$2 6 1 4 9 10 example_config_freepdk45_and2_dec
* cell instance $8 r0 *1 0.56,0
X$8 1 3 9 10 example_config_freepdk45_pinv
* cell instance $9 r0 *1 2.0875,2.73
X$9 7 3 2 9 10 example_config_freepdk45_and2_dec
* cell instance $15 m0 *1 0.56,2.73
X$15 2 4 9 10 example_config_freepdk45_pinv
* cell instance $16 r0 *1 2.0875,0
X$16 5 3 4 9 10 example_config_freepdk45_and2_dec
.ENDS example_config_freepdk45_hierarchical_predecode2x4

* cell write_driver
* pin din
* pin en
* pin br
* pin bl
* pin vdd
* pin gnd
.SUBCKT write_driver 1 2 5 9 11 12
* net 1 din
* net 2 en
* net 5 br
* net 9 bl
* net 11 vdd
* net 12 gnd
* device instance $1 r0 *1 0.17,3.0725 PMOS_VTG
M$1 11 3 8 11 PMOS_VTG L=0.05U W=0.36U AS=0.0378P AD=0.0252P PS=0.93U PD=0.5U
* device instance $2 r0 *1 0.36,3.0725 PMOS_VTG
M$2 8 4 9 11 PMOS_VTG L=0.05U W=0.36U AS=0.0252P AD=0.0378P PS=0.5U PD=0.93U
* device instance $3 r0 *1 0.17,2.46 PMOS_VTG
M$3 11 1 7 11 PMOS_VTG L=0.05U W=0.36U AS=0.0378P AD=0.0252P PS=0.93U PD=0.5U
* device instance $4 r0 *1 0.36,2.46 PMOS_VTG
M$4 7 4 5 11 PMOS_VTG L=0.05U W=0.36U AS=0.0252P AD=0.0378P PS=0.5U PD=0.93U
* device instance $5 r0 *1 0.51,0.885 PMOS_VTG
M$5 4 2 11 11 PMOS_VTG L=0.05U W=0.36U AS=0.0378P AD=0.0378P PS=0.93U PD=0.93U
* device instance $6 r0 *1 0.17,0.885 PMOS_VTG
M$6 11 1 3 11 PMOS_VTG L=0.05U W=0.36U AS=0.0378P AD=0.0378P PS=0.93U PD=0.93U
* device instance $7 r0 *1 0.17,3.6775 NMOS_VTG
M$7 12 3 10 12 NMOS_VTG L=0.05U W=0.18U AS=0.0189P AD=0.0126P PS=0.57U PD=0.32U
* device instance $8 r0 *1 0.36,3.6775 NMOS_VTG
M$8 10 2 9 12 NMOS_VTG L=0.05U W=0.18U AS=0.0126P AD=0.0189P PS=0.32U PD=0.57U
* device instance $9 r0 *1 0.17,1.855 NMOS_VTG
M$9 12 1 6 12 NMOS_VTG L=0.05U W=0.18U AS=0.0189P AD=0.0126P PS=0.57U PD=0.32U
* device instance $10 r0 *1 0.36,1.855 NMOS_VTG
M$10 6 2 5 12 NMOS_VTG L=0.05U W=0.18U AS=0.0126P AD=0.0189P PS=0.32U PD=0.57U
* device instance $11 r0 *1 0.51,1.49 NMOS_VTG
M$11 4 2 12 12 NMOS_VTG L=0.05U W=0.18U AS=0.0189P AD=0.0189P PS=0.57U PD=0.57U
* device instance $12 r0 *1 0.17,1.49 NMOS_VTG
M$12 12 1 3 12 NMOS_VTG L=0.05U W=0.18U AS=0.0189P AD=0.0189P PS=0.57U PD=0.57U
.ENDS write_driver

* cell sense_amp
* pin br
* pin dout
* pin bl
* pin en
* pin vdd
* pin gnd
.SUBCKT sense_amp 1 3 4 6 9 10
* net 1 br
* net 3 dout
* net 4 bl
* net 6 en
* net 9 vdd
* net 10 gnd
* device instance $1 r0 *1 0.2575,4.0975 PMOS_VTG
M$1 5 7 9 9 PMOS_VTG L=0.05U W=0.54U AS=0.0567P AD=0.0378P PS=1.29U PD=0.68U
* device instance $2 r0 *1 0.4475,4.0975 PMOS_VTG
M$2 9 5 7 9 PMOS_VTG L=0.05U W=0.54U AS=0.0378P AD=0.0567P PS=0.68U PD=1.29U
* device instance $3 r0 *1 0.4475,3.15 PMOS_VTG
M$3 7 6 1 9 PMOS_VTG L=0.05U W=0.72U AS=0.0756P AD=0.0756P PS=1.65U PD=1.65U
* device instance $4 r0 *1 0.2575,2.18 PMOS_VTG
M$4 4 6 5 9 PMOS_VTG L=0.05U W=0.72U AS=0.0756P AD=0.0756P PS=1.65U PD=1.65U
* device instance $5 r0 *1 0.4625,0.955 PMOS_VTG
M$5 9 5 2 9 PMOS_VTG L=0.05U W=0.18U AS=0.03285P AD=0.0189P PS=0.695U PD=0.57U
* device instance $6 r0 *1 0.2575,1.135 PMOS_VTG
M$6 3 2 9 9 PMOS_VTG L=0.05U W=0.54U AS=0.0567P AD=0.03285P PS=1.29U PD=0.695U
* device instance $7 r0 *1 0.3575,5.445 NMOS_VTG
M$7 8 6 10 10 NMOS_VTG L=0.05U W=0.27U AS=0.02835P AD=0.02835P PS=0.75U PD=0.75U
* device instance $8 r0 *1 0.2575,4.9875 NMOS_VTG
M$8 5 7 8 10 NMOS_VTG L=0.05U W=0.27U AS=0.02835P AD=0.0189P PS=0.75U PD=0.41U
* device instance $9 r0 *1 0.4475,4.9875 NMOS_VTG
M$9 8 5 7 10 NMOS_VTG L=0.05U W=0.27U AS=0.0189P AD=0.02835P PS=0.41U PD=0.75U
* device instance $10 r0 *1 0.2575,0.245 NMOS_VTG
M$10 3 2 10 10 NMOS_VTG L=0.05U W=0.27U AS=0.02835P AD=0.016425P PS=0.75U
+ PD=0.425U
* device instance $11 r0 *1 0.4625,0.335 NMOS_VTG
M$11 10 5 2 10 NMOS_VTG L=0.05U W=0.09U AS=0.016425P AD=0.00945P PS=0.425U
+ PD=0.39U
.ENDS sense_amp

* cell example_config_freepdk45_precharge_0
* pin en_bar
* pin bl
* pin br
* pin vdd
.SUBCKT example_config_freepdk45_precharge_0 1 2 3 4
* net 1 en_bar
* net 2 bl
* net 3 br
* net 4 vdd
* device instance $1 r0 *1 0.265,0.905 PMOS_VTG
M$1 2 1 4 4 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.022275P PS=0.795U
+ PD=0.435U
* device instance $2 r0 *1 0.48,0.905 PMOS_VTG
M$2 4 1 3 4 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.034425P PS=0.435U
+ PD=0.795U
* device instance $3 r0 *1 0.265,0.355 PMOS_VTG
M$3 2 1 3 4 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.034425P PS=0.795U
+ PD=0.795U
.ENDS example_config_freepdk45_precharge_0

* cell example_config_freepdk45_dummy_array
* pin wl_0_0
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_dummy_array 1 2 3
* net 1 wl_0_0
* net 2 vdd
* net 3 gnd
* cell instance $1 r0 *1 0.705,0
X$1 1 2 3 dummy_cell_1rw
* cell instance $2 r0 *1 0,0
X$2 1 2 3 dummy_cell_1rw
.ENDS example_config_freepdk45_dummy_array

* cell example_config_freepdk45_replica_column
* pin wl_0_0
* pin wl_0_1
* pin wl_0_2
* pin wl_0_3
* pin wl_0_4
* pin wl_0_5
* pin wl_0_6
* pin wl_0_7
* pin wl_0_8
* pin wl_0_9
* pin wl_0_10
* pin wl_0_11
* pin wl_0_12
* pin wl_0_13
* pin wl_0_14
* pin wl_0_15
* pin wl_0_16
* pin bl_0_0
* pin br_0_0
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_replica_column 1 2 3 4 5 6 7 8 9 10 11 12 13
+ 14 15 16 17 18 19 20 21
* net 1 wl_0_0
* net 2 wl_0_1
* net 3 wl_0_2
* net 4 wl_0_3
* net 5 wl_0_4
* net 6 wl_0_5
* net 7 wl_0_6
* net 8 wl_0_7
* net 9 wl_0_8
* net 10 wl_0_9
* net 11 wl_0_10
* net 12 wl_0_11
* net 13 wl_0_12
* net 14 wl_0_13
* net 15 wl_0_14
* net 16 wl_0_15
* net 17 wl_0_16
* net 18 bl_0_0
* net 19 br_0_0
* net 20 vdd
* net 21 gnd
* cell instance $1 m0 *1 0,1.365
X$1 18 1 19 20 21 replica_cell_1rw
* cell instance $2 r0 *1 0,1.365
X$2 18 2 19 20 21 replica_cell_1rw
* cell instance $3 m0 *1 0,4.095
X$3 18 3 19 20 21 replica_cell_1rw
* cell instance $4 r0 *1 0,4.095
X$4 18 4 19 20 21 replica_cell_1rw
* cell instance $5 m0 *1 0,6.825
X$5 18 5 19 20 21 replica_cell_1rw
* cell instance $6 r0 *1 0,6.825
X$6 18 6 19 20 21 replica_cell_1rw
* cell instance $7 m0 *1 0,9.555
X$7 18 7 19 20 21 replica_cell_1rw
* cell instance $8 r0 *1 0,9.555
X$8 18 8 19 20 21 replica_cell_1rw
* cell instance $9 m0 *1 0,12.285
X$9 18 9 19 20 21 replica_cell_1rw
* cell instance $10 r0 *1 0,12.285
X$10 18 10 19 20 21 replica_cell_1rw
* cell instance $11 m0 *1 0,15.015
X$11 18 11 19 20 21 replica_cell_1rw
* cell instance $12 r0 *1 0,15.015
X$12 18 12 19 20 21 replica_cell_1rw
* cell instance $13 m0 *1 0,17.745
X$13 18 13 19 20 21 replica_cell_1rw
* cell instance $14 r0 *1 0,17.745
X$14 18 14 19 20 21 replica_cell_1rw
* cell instance $15 m0 *1 0,20.475
X$15 18 15 19 20 21 replica_cell_1rw
* cell instance $16 r0 *1 0,20.475
X$16 18 16 19 20 21 replica_cell_1rw
* cell instance $17 m0 *1 0,23.205
X$17 18 17 19 20 21 replica_cell_1rw
.ENDS example_config_freepdk45_replica_column

* cell example_config_freepdk45_bitcell_array
* pin wl_0_0
* pin wl_0_1
* pin wl_0_2
* pin wl_0_3
* pin wl_0_4
* pin wl_0_5
* pin wl_0_6
* pin wl_0_7
* pin bl_0_0
* pin br_0_0
* pin bl_0_1
* pin br_0_1
* pin wl_0_8
* pin wl_0_9
* pin wl_0_10
* pin wl_0_11
* pin wl_0_12
* pin wl_0_13
* pin wl_0_14
* pin wl_0_15
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_bitcell_array 1 2 3 4 5 6 7 8 9 10 11 12 13 14
+ 15 16 17 18 19 20 21 22
* net 1 wl_0_0
* net 2 wl_0_1
* net 3 wl_0_2
* net 4 wl_0_3
* net 5 wl_0_4
* net 6 wl_0_5
* net 7 wl_0_6
* net 8 wl_0_7
* net 9 bl_0_0
* net 10 br_0_0
* net 11 bl_0_1
* net 12 br_0_1
* net 13 wl_0_8
* net 14 wl_0_9
* net 15 wl_0_10
* net 16 wl_0_11
* net 17 wl_0_12
* net 18 wl_0_13
* net 19 wl_0_14
* net 20 wl_0_15
* net 21 vdd
* net 22 gnd
* cell instance $1 r0 *1 0.705,0
X$1 11 1 12 21 22 cell_1rw
* cell instance $2 r0 *1 0,0
X$2 9 1 10 21 22 cell_1rw
* cell instance $3 m0 *1 0,2.73
X$3 9 2 10 21 22 cell_1rw
* cell instance $4 m0 *1 0.705,2.73
X$4 11 2 12 21 22 cell_1rw
* cell instance $5 r0 *1 0,2.73
X$5 9 3 10 21 22 cell_1rw
* cell instance $6 r0 *1 0.705,2.73
X$6 11 3 12 21 22 cell_1rw
* cell instance $7 m0 *1 0,5.46
X$7 9 4 10 21 22 cell_1rw
* cell instance $8 m0 *1 0.705,5.46
X$8 11 4 12 21 22 cell_1rw
* cell instance $9 r0 *1 0,5.46
X$9 9 5 10 21 22 cell_1rw
* cell instance $10 r0 *1 0.705,5.46
X$10 11 5 12 21 22 cell_1rw
* cell instance $11 m0 *1 0,8.19
X$11 9 6 10 21 22 cell_1rw
* cell instance $12 m0 *1 0.705,8.19
X$12 11 6 12 21 22 cell_1rw
* cell instance $13 r0 *1 0,8.19
X$13 9 7 10 21 22 cell_1rw
* cell instance $14 r0 *1 0.705,8.19
X$14 11 7 12 21 22 cell_1rw
* cell instance $15 m0 *1 0,10.92
X$15 9 8 10 21 22 cell_1rw
* cell instance $16 m0 *1 0.705,10.92
X$16 11 8 12 21 22 cell_1rw
* cell instance $17 r0 *1 0,10.92
X$17 9 13 10 21 22 cell_1rw
* cell instance $18 m0 *1 0,13.65
X$18 9 14 10 21 22 cell_1rw
* cell instance $19 r0 *1 0,13.65
X$19 9 15 10 21 22 cell_1rw
* cell instance $20 m0 *1 0,16.38
X$20 9 16 10 21 22 cell_1rw
* cell instance $21 r0 *1 0,16.38
X$21 9 17 10 21 22 cell_1rw
* cell instance $22 m0 *1 0,19.11
X$22 9 18 10 21 22 cell_1rw
* cell instance $23 r0 *1 0,19.11
X$23 9 19 10 21 22 cell_1rw
* cell instance $24 m0 *1 0,21.84
X$24 9 20 10 21 22 cell_1rw
* cell instance $25 r0 *1 0.705,10.92
X$25 11 13 12 21 22 cell_1rw
* cell instance $26 m0 *1 0.705,13.65
X$26 11 14 12 21 22 cell_1rw
* cell instance $27 r0 *1 0.705,13.65
X$27 11 15 12 21 22 cell_1rw
* cell instance $28 m0 *1 0.705,16.38
X$28 11 16 12 21 22 cell_1rw
* cell instance $29 r0 *1 0.705,16.38
X$29 11 17 12 21 22 cell_1rw
* cell instance $30 m0 *1 0.705,19.11
X$30 11 18 12 21 22 cell_1rw
* cell instance $31 r0 *1 0.705,19.11
X$31 11 19 12 21 22 cell_1rw
* cell instance $32 m0 *1 0.705,21.84
X$32 11 20 12 21 22 cell_1rw
.ENDS example_config_freepdk45_bitcell_array

* cell example_config_freepdk45_and2_dec
* pin Z
* pin A
* pin B
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_and2_dec 2 3 4 5 6
* net 2 Z
* net 3 A
* net 4 B
* net 5 vdd
* net 6 gnd
* cell instance $1 r0 *1 0,0
X$1 3 4 1 5 6 example_config_freepdk45_pnand2
* cell instance $2 r0 *1 0.9025,0
X$2 1 2 5 6 example_config_freepdk45_pinv
.ENDS example_config_freepdk45_and2_dec

* cell dummy_cell_1rw
* pin wl
* pin vdd
* pin gnd
.SUBCKT dummy_cell_1rw 2 6 7
* net 2 wl
* net 6 vdd
* net 7 gnd
* device instance $1 r0 *1 0.61,1.2075 PMOS_VTG
M$1 5 1 6 6 PMOS_VTG L=0.05U W=0.09U AS=0.00945P AD=0.00945P PS=0.39U PD=0.39U
* device instance $2 r0 *1 0.095,1.2075 PMOS_VTG
M$2 6 5 1 6 PMOS_VTG L=0.05U W=0.09U AS=0.00945P AD=0.00945P PS=0.39U PD=0.39U
* device instance $3 r0 *1 0.61,0.67 NMOS_VTG
M$3 5 1 7 7 NMOS_VTG L=0.05U W=0.205U AS=0.021525P AD=0.021525P PS=0.62U
+ PD=0.62U
* device instance $4 r0 *1 0.095,0.67 NMOS_VTG
M$4 7 5 1 7 NMOS_VTG L=0.05U W=0.205U AS=0.021525P AD=0.021525P PS=0.62U
+ PD=0.62U
* device instance $5 r0 *1 0.53,0.315 NMOS_VTG
M$5 3 2 5 7 NMOS_VTG L=0.05U W=0.135U AS=0.014175P AD=0.014175P PS=0.48U
+ PD=0.48U
* device instance $6 r0 *1 0.175,0.315 NMOS_VTG
M$6 1 2 4 7 NMOS_VTG L=0.05U W=0.135U AS=0.014175P AD=0.014175P PS=0.48U
+ PD=0.48U
.ENDS dummy_cell_1rw

* cell replica_cell_1rw
* pin bl
* pin wl
* pin br
* pin vdd
* pin gnd
.SUBCKT replica_cell_1rw 1 2 4 5 6
* net 1 bl
* net 2 wl
* net 4 br
* net 5 vdd
* net 6 gnd
* device instance $1 r0 *1 0.61,1.2075 PMOS_VTG
M$1 5 3 5 5 PMOS_VTG L=0.05U W=0.09U AS=0.00945P AD=0.0099P PS=0.39U PD=0.4U
* device instance $2 r0 *1 0.095,1.2075 PMOS_VTG
M$2 5 5 3 5 PMOS_VTG L=0.05U W=0.09U AS=0.0099P AD=0.00945P PS=0.4U PD=0.39U
* device instance $3 r0 *1 0.61,0.67 NMOS_VTG
M$3 5 3 6 6 NMOS_VTG L=0.05U W=0.205U AS=0.021525P AD=0.02255P PS=0.62U PD=0.63U
* device instance $4 r0 *1 0.095,0.67 NMOS_VTG
M$4 6 5 3 6 NMOS_VTG L=0.05U W=0.205U AS=0.02255P AD=0.021525P PS=0.63U PD=0.62U
* device instance $5 r0 *1 0.53,0.315 NMOS_VTG
M$5 4 2 5 6 NMOS_VTG L=0.05U W=0.135U AS=0.014175P AD=0.014175P PS=0.48U
+ PD=0.48U
* device instance $6 r0 *1 0.175,0.315 NMOS_VTG
M$6 3 2 1 6 NMOS_VTG L=0.05U W=0.135U AS=0.014175P AD=0.014175P PS=0.48U
+ PD=0.48U
.ENDS replica_cell_1rw

* cell cell_1rw
* pin bl
* pin wl
* pin br
* pin vdd
* pin gnd
.SUBCKT cell_1rw 1 2 4 6 7
* net 1 bl
* net 2 wl
* net 3 Q
* net 4 br
* net 5 Q_bar
* net 6 vdd
* net 7 gnd
* device instance $1 r0 *1 0.61,1.2075 PMOS_VTG
M$1 5 3 6 6 PMOS_VTG L=0.05U W=0.09U AS=0.00945P AD=0.0099P PS=0.39U PD=0.4U
* device instance $2 r0 *1 0.095,1.2075 PMOS_VTG
M$2 6 5 3 6 PMOS_VTG L=0.05U W=0.09U AS=0.0099P AD=0.00945P PS=0.4U PD=0.39U
* device instance $3 r0 *1 0.61,0.67 NMOS_VTG
M$3 5 3 7 7 NMOS_VTG L=0.05U W=0.205U AS=0.021525P AD=0.02255P PS=0.62U PD=0.63U
* device instance $4 r0 *1 0.095,0.67 NMOS_VTG
M$4 7 5 3 7 NMOS_VTG L=0.05U W=0.205U AS=0.02255P AD=0.021525P PS=0.63U PD=0.62U
* device instance $5 r0 *1 0.53,0.315 NMOS_VTG
M$5 4 2 5 7 NMOS_VTG L=0.05U W=0.135U AS=0.014175P AD=0.014175P PS=0.48U
+ PD=0.48U
* device instance $6 r0 *1 0.175,0.315 NMOS_VTG
M$6 3 2 1 7 NMOS_VTG L=0.05U W=0.135U AS=0.014175P AD=0.014175P PS=0.48U
+ PD=0.48U
.ENDS cell_1rw

* cell example_config_freepdk45_pnand2
* pin A
* pin B
* pin Z
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pnand2 1 2 3 4 5
* net 1 A
* net 2 B
* net 3 Z
* net 4 vdd
* net 5 gnd
* device instance $1 r0 *1 0.2325,1.105 PMOS_VTG
M$1 4 1 3 4 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.022275P PS=0.795U
+ PD=0.435U
* device instance $2 r0 *1 0.4475,1.105 PMOS_VTG
M$2 3 2 4 4 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.034425P PS=0.435U
+ PD=0.795U
* device instance $3 r0 *1 0.2325,0.215 NMOS_VTG
M$3 5 1 6 5 NMOS_VTG L=0.05U W=0.18U AS=0.02295P AD=0.01485P PS=0.615U PD=0.345U
* device instance $4 r0 *1 0.4475,0.215 NMOS_VTG
M$4 6 2 3 5 NMOS_VTG L=0.05U W=0.18U AS=0.01485P AD=0.02295P PS=0.345U PD=0.615U
.ENDS example_config_freepdk45_pnand2

* cell example_config_freepdk45_pinv
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT example_config_freepdk45_pinv 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.17 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.09U AS=0.011475P AD=0.011475P PS=0.435U
+ PD=0.435U
* device instance $2 r0 *1 0.2325,1.105 PMOS_VTG
M$2 3 1 2 3 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.034425P PS=0.795U
+ PD=0.795U
.ENDS example_config_freepdk45_pinv
