VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_1rw0r0w_32_512_freepdk45
   CLASS BLOCK ;
   SIZE 139.57 BY 203.195 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  31.1175 0.0 31.2575 0.14 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  33.9775 0.0 34.1175 0.14 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  36.8375 0.0 36.9775 0.14 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  39.6975 0.0 39.8375 0.14 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  42.5575 0.0 42.6975 0.14 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  45.4175 0.0 45.5575 0.14 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  48.2775 0.0 48.4175 0.14 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  51.1375 0.0 51.2775 0.14 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  53.9975 0.0 54.1375 0.14 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  56.8575 0.0 56.9975 0.14 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  59.7175 0.0 59.8575 0.14 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  62.5775 0.0 62.7175 0.14 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  65.4375 0.0 65.5775 0.14 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  68.2975 0.0 68.4375 0.14 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  71.1575 0.0 71.2975 0.14 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  74.0175 0.0 74.1575 0.14 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  76.8775 0.0 77.0175 0.14 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  79.7375 0.0 79.8775 0.14 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  82.5975 0.0 82.7375 0.14 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  85.4575 0.0 85.5975 0.14 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  88.3175 0.0 88.4575 0.14 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  91.1775 0.0 91.3175 0.14 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  94.0375 0.0 94.1775 0.14 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  96.8975 0.0 97.0375 0.14 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  99.7575 0.0 99.8975 0.14 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  102.6175 0.0 102.7575 0.14 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  105.4775 0.0 105.6175 0.14 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  108.3375 0.0 108.4775 0.14 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  111.1975 0.0 111.3375 0.14 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  114.0575 0.0 114.1975 0.14 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  116.9175 0.0 117.0575 0.14 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  119.7775 0.0 119.9175 0.14 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  25.3975 0.0 25.5375 0.14 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  28.2575 0.0 28.3975 0.14 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 55.18 0.14 55.32 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 57.91 0.14 58.05 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 60.12 0.14 60.26 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 62.85 0.14 62.99 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 65.06 0.14 65.2 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 67.79 0.14 67.93 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 70.0 0.14 70.14 ;
      END
   END addr0[8]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 5.0 0.14 5.14 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 7.73 0.14 7.87 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  9.84 0.0 9.98 0.14 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  44.3725 0.0 44.5125 0.14 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  47.1925 0.0 47.3325 0.14 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  50.0125 0.0 50.1525 0.14 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  52.8325 0.0 52.9725 0.14 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  55.6525 0.0 55.7925 0.14 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  58.4725 0.0 58.6125 0.14 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  61.2925 0.0 61.4325 0.14 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  64.1125 0.0 64.2525 0.14 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  66.9325 0.0 67.0725 0.14 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  69.7525 0.0 69.8925 0.14 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  72.5725 0.0 72.7125 0.14 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  75.3925 0.0 75.5325 0.14 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  78.2125 0.0 78.3525 0.14 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  81.0325 0.0 81.1725 0.14 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  83.8525 0.0 83.9925 0.14 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  86.6725 0.0 86.8125 0.14 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  89.4925 0.0 89.6325 0.14 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  92.3125 0.0 92.4525 0.14 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  95.1325 0.0 95.2725 0.14 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  97.9525 0.0 98.0925 0.14 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  100.7725 0.0 100.9125 0.14 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  103.5925 0.0 103.7325 0.14 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  106.4125 0.0 106.5525 0.14 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  109.2325 0.0 109.3725 0.14 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  112.0525 0.0 112.1925 0.14 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  114.8725 0.0 115.0125 0.14 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  117.6925 0.0 117.8325 0.14 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  120.5125 0.0 120.6525 0.14 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  123.3325 0.0 123.4725 0.14 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  126.1525 0.0 126.2925 0.14 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  139.43 13.1625 139.57 13.3025 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  139.43 12.9275 139.57 13.0675 ;
      END
   END dout0[31]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 139.43 203.055 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 139.43 203.055 ;
   LAYER  metal3 ;
      RECT  0.28 55.04 139.43 55.46 ;
      RECT  0.28 55.46 139.43 203.055 ;
      RECT  0.14 55.46 0.28 57.77 ;
      RECT  0.14 58.19 0.28 59.98 ;
      RECT  0.14 60.4 0.28 62.71 ;
      RECT  0.14 63.13 0.28 64.92 ;
      RECT  0.14 65.34 0.28 67.65 ;
      RECT  0.14 68.07 0.28 69.86 ;
      RECT  0.14 70.28 0.28 203.055 ;
      RECT  0.14 0.14 0.28 4.86 ;
      RECT  0.14 5.28 0.28 7.59 ;
      RECT  0.14 8.01 0.28 55.04 ;
      RECT  0.28 0.14 139.29 13.0225 ;
      RECT  0.28 13.0225 139.29 13.4425 ;
      RECT  0.28 13.4425 139.29 55.04 ;
      RECT  139.29 13.4425 139.43 55.04 ;
      RECT  139.29 0.14 139.43 12.7875 ;
   LAYER  metal4 ;
      RECT  0.14 0.42 30.8375 203.055 ;
      RECT  30.8375 0.42 31.5375 203.055 ;
      RECT  31.5375 0.42 139.43 203.055 ;
      RECT  31.5375 0.14 33.6975 0.42 ;
      RECT  34.3975 0.14 36.5575 0.42 ;
      RECT  37.2575 0.14 39.4175 0.42 ;
      RECT  40.1175 0.14 42.2775 0.42 ;
      RECT  25.8175 0.14 27.9775 0.42 ;
      RECT  28.6775 0.14 30.8375 0.42 ;
      RECT  0.14 0.14 9.56 0.42 ;
      RECT  10.26 0.14 25.1175 0.42 ;
      RECT  42.9775 0.14 44.0925 0.42 ;
      RECT  44.7925 0.14 45.1375 0.42 ;
      RECT  45.8375 0.14 46.9125 0.42 ;
      RECT  47.6125 0.14 47.9975 0.42 ;
      RECT  48.6975 0.14 49.7325 0.42 ;
      RECT  50.4325 0.14 50.8575 0.42 ;
      RECT  51.5575 0.14 52.5525 0.42 ;
      RECT  53.2525 0.14 53.7175 0.42 ;
      RECT  54.4175 0.14 55.3725 0.42 ;
      RECT  56.0725 0.14 56.5775 0.42 ;
      RECT  57.2775 0.14 58.1925 0.42 ;
      RECT  58.8925 0.14 59.4375 0.42 ;
      RECT  60.1375 0.14 61.0125 0.42 ;
      RECT  61.7125 0.14 62.2975 0.42 ;
      RECT  62.9975 0.14 63.8325 0.42 ;
      RECT  64.5325 0.14 65.1575 0.42 ;
      RECT  65.8575 0.14 66.6525 0.42 ;
      RECT  67.3525 0.14 68.0175 0.42 ;
      RECT  68.7175 0.14 69.4725 0.42 ;
      RECT  70.1725 0.14 70.8775 0.42 ;
      RECT  71.5775 0.14 72.2925 0.42 ;
      RECT  72.9925 0.14 73.7375 0.42 ;
      RECT  74.4375 0.14 75.1125 0.42 ;
      RECT  75.8125 0.14 76.5975 0.42 ;
      RECT  77.2975 0.14 77.9325 0.42 ;
      RECT  78.6325 0.14 79.4575 0.42 ;
      RECT  80.1575 0.14 80.7525 0.42 ;
      RECT  81.4525 0.14 82.3175 0.42 ;
      RECT  83.0175 0.14 83.5725 0.42 ;
      RECT  84.2725 0.14 85.1775 0.42 ;
      RECT  85.8775 0.14 86.3925 0.42 ;
      RECT  87.0925 0.14 88.0375 0.42 ;
      RECT  88.7375 0.14 89.2125 0.42 ;
      RECT  89.9125 0.14 90.8975 0.42 ;
      RECT  91.5975 0.14 92.0325 0.42 ;
      RECT  92.7325 0.14 93.7575 0.42 ;
      RECT  94.4575 0.14 94.8525 0.42 ;
      RECT  95.5525 0.14 96.6175 0.42 ;
      RECT  97.3175 0.14 97.6725 0.42 ;
      RECT  98.3725 0.14 99.4775 0.42 ;
      RECT  100.1775 0.14 100.4925 0.42 ;
      RECT  101.1925 0.14 102.3375 0.42 ;
      RECT  103.0375 0.14 103.3125 0.42 ;
      RECT  104.0125 0.14 105.1975 0.42 ;
      RECT  105.8975 0.14 106.1325 0.42 ;
      RECT  106.8325 0.14 108.0575 0.42 ;
      RECT  108.7575 0.14 108.9525 0.42 ;
      RECT  109.6525 0.14 110.9175 0.42 ;
      RECT  111.6175 0.14 111.7725 0.42 ;
      RECT  112.4725 0.14 113.7775 0.42 ;
      RECT  114.4775 0.14 114.5925 0.42 ;
      RECT  115.2925 0.14 116.6375 0.42 ;
      RECT  117.3375 0.14 117.4125 0.42 ;
      RECT  118.1125 0.14 119.4975 0.42 ;
      RECT  120.1975 0.14 120.2325 0.42 ;
      RECT  120.9325 0.14 123.0525 0.42 ;
      RECT  123.7525 0.14 125.8725 0.42 ;
      RECT  126.5725 0.14 139.43 0.42 ;
   END
END    sram_1rw0r0w_32_512_freepdk45
END    LIBRARY
