VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_0rw1r1w_576_16_freepdk45
   CLASS BLOCK ;
   SIZE 1785.29 BY 192.97 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  138.1425 0.0 138.2825 0.14 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  141.0025 0.0 141.1425 0.14 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  143.8625 0.0 144.0025 0.14 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  146.7225 0.0 146.8625 0.14 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  149.5825 0.0 149.7225 0.14 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  152.4425 0.0 152.5825 0.14 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  155.3025 0.0 155.4425 0.14 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  158.1625 0.0 158.3025 0.14 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  161.0225 0.0 161.1625 0.14 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  163.8825 0.0 164.0225 0.14 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  166.7425 0.0 166.8825 0.14 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  169.6025 0.0 169.7425 0.14 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  172.4625 0.0 172.6025 0.14 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  175.3225 0.0 175.4625 0.14 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  178.1825 0.0 178.3225 0.14 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  181.0425 0.0 181.1825 0.14 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  183.9025 0.0 184.0425 0.14 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  186.7625 0.0 186.9025 0.14 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  189.6225 0.0 189.7625 0.14 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  192.4825 0.0 192.6225 0.14 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  195.3425 0.0 195.4825 0.14 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  198.2025 0.0 198.3425 0.14 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  201.0625 0.0 201.2025 0.14 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  203.9225 0.0 204.0625 0.14 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  206.7825 0.0 206.9225 0.14 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  209.6425 0.0 209.7825 0.14 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  212.5025 0.0 212.6425 0.14 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  215.3625 0.0 215.5025 0.14 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  218.2225 0.0 218.3625 0.14 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  221.0825 0.0 221.2225 0.14 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  223.9425 0.0 224.0825 0.14 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  226.8025 0.0 226.9425 0.14 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  229.6625 0.0 229.8025 0.14 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  232.5225 0.0 232.6625 0.14 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  235.3825 0.0 235.5225 0.14 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  238.2425 0.0 238.3825 0.14 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  241.1025 0.0 241.2425 0.14 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  243.9625 0.0 244.1025 0.14 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  246.8225 0.0 246.9625 0.14 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  249.6825 0.0 249.8225 0.14 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  252.5425 0.0 252.6825 0.14 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  255.4025 0.0 255.5425 0.14 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  258.2625 0.0 258.4025 0.14 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  261.1225 0.0 261.2625 0.14 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  263.9825 0.0 264.1225 0.14 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  266.8425 0.0 266.9825 0.14 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  269.7025 0.0 269.8425 0.14 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  272.5625 0.0 272.7025 0.14 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  275.4225 0.0 275.5625 0.14 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  278.2825 0.0 278.4225 0.14 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  281.1425 0.0 281.2825 0.14 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  284.0025 0.0 284.1425 0.14 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  286.8625 0.0 287.0025 0.14 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  289.7225 0.0 289.8625 0.14 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  292.5825 0.0 292.7225 0.14 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  295.4425 0.0 295.5825 0.14 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  298.3025 0.0 298.4425 0.14 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  301.1625 0.0 301.3025 0.14 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  304.0225 0.0 304.1625 0.14 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  306.8825 0.0 307.0225 0.14 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  309.7425 0.0 309.8825 0.14 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  312.6025 0.0 312.7425 0.14 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  315.4625 0.0 315.6025 0.14 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  318.3225 0.0 318.4625 0.14 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  321.1825 0.0 321.3225 0.14 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  324.0425 0.0 324.1825 0.14 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  326.9025 0.0 327.0425 0.14 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  329.7625 0.0 329.9025 0.14 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  332.6225 0.0 332.7625 0.14 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  335.4825 0.0 335.6225 0.14 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  338.3425 0.0 338.4825 0.14 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  341.2025 0.0 341.3425 0.14 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  344.0625 0.0 344.2025 0.14 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  346.9225 0.0 347.0625 0.14 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  349.7825 0.0 349.9225 0.14 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  352.6425 0.0 352.7825 0.14 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  355.5025 0.0 355.6425 0.14 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  358.3625 0.0 358.5025 0.14 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  361.2225 0.0 361.3625 0.14 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  364.0825 0.0 364.2225 0.14 ;
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  366.9425 0.0 367.0825 0.14 ;
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  369.8025 0.0 369.9425 0.14 ;
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  372.6625 0.0 372.8025 0.14 ;
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  375.5225 0.0 375.6625 0.14 ;
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  378.3825 0.0 378.5225 0.14 ;
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  381.2425 0.0 381.3825 0.14 ;
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  384.1025 0.0 384.2425 0.14 ;
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  386.9625 0.0 387.1025 0.14 ;
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  389.8225 0.0 389.9625 0.14 ;
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  392.6825 0.0 392.8225 0.14 ;
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  395.5425 0.0 395.6825 0.14 ;
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  398.4025 0.0 398.5425 0.14 ;
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  401.2625 0.0 401.4025 0.14 ;
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  404.1225 0.0 404.2625 0.14 ;
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  406.9825 0.0 407.1225 0.14 ;
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  409.8425 0.0 409.9825 0.14 ;
      END
   END din0[95]
   PIN din0[96]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  412.7025 0.0 412.8425 0.14 ;
      END
   END din0[96]
   PIN din0[97]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  415.5625 0.0 415.7025 0.14 ;
      END
   END din0[97]
   PIN din0[98]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  418.4225 0.0 418.5625 0.14 ;
      END
   END din0[98]
   PIN din0[99]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  421.2825 0.0 421.4225 0.14 ;
      END
   END din0[99]
   PIN din0[100]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  424.1425 0.0 424.2825 0.14 ;
      END
   END din0[100]
   PIN din0[101]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  427.0025 0.0 427.1425 0.14 ;
      END
   END din0[101]
   PIN din0[102]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  429.8625 0.0 430.0025 0.14 ;
      END
   END din0[102]
   PIN din0[103]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  432.7225 0.0 432.8625 0.14 ;
      END
   END din0[103]
   PIN din0[104]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  435.5825 0.0 435.7225 0.14 ;
      END
   END din0[104]
   PIN din0[105]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  438.4425 0.0 438.5825 0.14 ;
      END
   END din0[105]
   PIN din0[106]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  441.3025 0.0 441.4425 0.14 ;
      END
   END din0[106]
   PIN din0[107]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  444.1625 0.0 444.3025 0.14 ;
      END
   END din0[107]
   PIN din0[108]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  447.0225 0.0 447.1625 0.14 ;
      END
   END din0[108]
   PIN din0[109]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  449.8825 0.0 450.0225 0.14 ;
      END
   END din0[109]
   PIN din0[110]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  452.7425 0.0 452.8825 0.14 ;
      END
   END din0[110]
   PIN din0[111]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  455.6025 0.0 455.7425 0.14 ;
      END
   END din0[111]
   PIN din0[112]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  458.4625 0.0 458.6025 0.14 ;
      END
   END din0[112]
   PIN din0[113]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  461.3225 0.0 461.4625 0.14 ;
      END
   END din0[113]
   PIN din0[114]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  464.1825 0.0 464.3225 0.14 ;
      END
   END din0[114]
   PIN din0[115]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  467.0425 0.0 467.1825 0.14 ;
      END
   END din0[115]
   PIN din0[116]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  469.9025 0.0 470.0425 0.14 ;
      END
   END din0[116]
   PIN din0[117]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  472.7625 0.0 472.9025 0.14 ;
      END
   END din0[117]
   PIN din0[118]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  475.6225 0.0 475.7625 0.14 ;
      END
   END din0[118]
   PIN din0[119]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  478.4825 0.0 478.6225 0.14 ;
      END
   END din0[119]
   PIN din0[120]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  481.3425 0.0 481.4825 0.14 ;
      END
   END din0[120]
   PIN din0[121]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  484.2025 0.0 484.3425 0.14 ;
      END
   END din0[121]
   PIN din0[122]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  487.0625 0.0 487.2025 0.14 ;
      END
   END din0[122]
   PIN din0[123]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  489.9225 0.0 490.0625 0.14 ;
      END
   END din0[123]
   PIN din0[124]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  492.7825 0.0 492.9225 0.14 ;
      END
   END din0[124]
   PIN din0[125]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  495.6425 0.0 495.7825 0.14 ;
      END
   END din0[125]
   PIN din0[126]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  498.5025 0.0 498.6425 0.14 ;
      END
   END din0[126]
   PIN din0[127]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  501.3625 0.0 501.5025 0.14 ;
      END
   END din0[127]
   PIN din0[128]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  504.2225 0.0 504.3625 0.14 ;
      END
   END din0[128]
   PIN din0[129]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  507.0825 0.0 507.2225 0.14 ;
      END
   END din0[129]
   PIN din0[130]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  509.9425 0.0 510.0825 0.14 ;
      END
   END din0[130]
   PIN din0[131]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  512.8025 0.0 512.9425 0.14 ;
      END
   END din0[131]
   PIN din0[132]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  515.6625 0.0 515.8025 0.14 ;
      END
   END din0[132]
   PIN din0[133]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  518.5225 0.0 518.6625 0.14 ;
      END
   END din0[133]
   PIN din0[134]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  521.3825 0.0 521.5225 0.14 ;
      END
   END din0[134]
   PIN din0[135]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  524.2425 0.0 524.3825 0.14 ;
      END
   END din0[135]
   PIN din0[136]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  527.1025 0.0 527.2425 0.14 ;
      END
   END din0[136]
   PIN din0[137]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  529.9625 0.0 530.1025 0.14 ;
      END
   END din0[137]
   PIN din0[138]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  532.8225 0.0 532.9625 0.14 ;
      END
   END din0[138]
   PIN din0[139]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  535.6825 0.0 535.8225 0.14 ;
      END
   END din0[139]
   PIN din0[140]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  538.5425 0.0 538.6825 0.14 ;
      END
   END din0[140]
   PIN din0[141]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  541.4025 0.0 541.5425 0.14 ;
      END
   END din0[141]
   PIN din0[142]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  544.2625 0.0 544.4025 0.14 ;
      END
   END din0[142]
   PIN din0[143]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  547.1225 0.0 547.2625 0.14 ;
      END
   END din0[143]
   PIN din0[144]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  549.9825 0.0 550.1225 0.14 ;
      END
   END din0[144]
   PIN din0[145]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  552.8425 0.0 552.9825 0.14 ;
      END
   END din0[145]
   PIN din0[146]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  555.7025 0.0 555.8425 0.14 ;
      END
   END din0[146]
   PIN din0[147]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  558.5625 0.0 558.7025 0.14 ;
      END
   END din0[147]
   PIN din0[148]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  561.4225 0.0 561.5625 0.14 ;
      END
   END din0[148]
   PIN din0[149]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  564.2825 0.0 564.4225 0.14 ;
      END
   END din0[149]
   PIN din0[150]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  567.1425 0.0 567.2825 0.14 ;
      END
   END din0[150]
   PIN din0[151]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  570.0025 0.0 570.1425 0.14 ;
      END
   END din0[151]
   PIN din0[152]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  572.8625 0.0 573.0025 0.14 ;
      END
   END din0[152]
   PIN din0[153]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  575.7225 0.0 575.8625 0.14 ;
      END
   END din0[153]
   PIN din0[154]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  578.5825 0.0 578.7225 0.14 ;
      END
   END din0[154]
   PIN din0[155]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  581.4425 0.0 581.5825 0.14 ;
      END
   END din0[155]
   PIN din0[156]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  584.3025 0.0 584.4425 0.14 ;
      END
   END din0[156]
   PIN din0[157]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  587.1625 0.0 587.3025 0.14 ;
      END
   END din0[157]
   PIN din0[158]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  590.0225 0.0 590.1625 0.14 ;
      END
   END din0[158]
   PIN din0[159]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  592.8825 0.0 593.0225 0.14 ;
      END
   END din0[159]
   PIN din0[160]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  595.7425 0.0 595.8825 0.14 ;
      END
   END din0[160]
   PIN din0[161]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  598.6025 0.0 598.7425 0.14 ;
      END
   END din0[161]
   PIN din0[162]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  601.4625 0.0 601.6025 0.14 ;
      END
   END din0[162]
   PIN din0[163]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  604.3225 0.0 604.4625 0.14 ;
      END
   END din0[163]
   PIN din0[164]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  607.1825 0.0 607.3225 0.14 ;
      END
   END din0[164]
   PIN din0[165]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  610.0425 0.0 610.1825 0.14 ;
      END
   END din0[165]
   PIN din0[166]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  612.9025 0.0 613.0425 0.14 ;
      END
   END din0[166]
   PIN din0[167]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  615.7625 0.0 615.9025 0.14 ;
      END
   END din0[167]
   PIN din0[168]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  618.6225 0.0 618.7625 0.14 ;
      END
   END din0[168]
   PIN din0[169]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  621.4825 0.0 621.6225 0.14 ;
      END
   END din0[169]
   PIN din0[170]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  624.3425 0.0 624.4825 0.14 ;
      END
   END din0[170]
   PIN din0[171]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  627.2025 0.0 627.3425 0.14 ;
      END
   END din0[171]
   PIN din0[172]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  630.0625 0.0 630.2025 0.14 ;
      END
   END din0[172]
   PIN din0[173]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  632.9225 0.0 633.0625 0.14 ;
      END
   END din0[173]
   PIN din0[174]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  635.7825 0.0 635.9225 0.14 ;
      END
   END din0[174]
   PIN din0[175]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  638.6425 0.0 638.7825 0.14 ;
      END
   END din0[175]
   PIN din0[176]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  641.5025 0.0 641.6425 0.14 ;
      END
   END din0[176]
   PIN din0[177]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  644.3625 0.0 644.5025 0.14 ;
      END
   END din0[177]
   PIN din0[178]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  647.2225 0.0 647.3625 0.14 ;
      END
   END din0[178]
   PIN din0[179]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  650.0825 0.0 650.2225 0.14 ;
      END
   END din0[179]
   PIN din0[180]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  652.9425 0.0 653.0825 0.14 ;
      END
   END din0[180]
   PIN din0[181]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  655.8025 0.0 655.9425 0.14 ;
      END
   END din0[181]
   PIN din0[182]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  658.6625 0.0 658.8025 0.14 ;
      END
   END din0[182]
   PIN din0[183]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  661.5225 0.0 661.6625 0.14 ;
      END
   END din0[183]
   PIN din0[184]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  664.3825 0.0 664.5225 0.14 ;
      END
   END din0[184]
   PIN din0[185]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  667.2425 0.0 667.3825 0.14 ;
      END
   END din0[185]
   PIN din0[186]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  670.1025 0.0 670.2425 0.14 ;
      END
   END din0[186]
   PIN din0[187]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  672.9625 0.0 673.1025 0.14 ;
      END
   END din0[187]
   PIN din0[188]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  675.8225 0.0 675.9625 0.14 ;
      END
   END din0[188]
   PIN din0[189]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  678.6825 0.0 678.8225 0.14 ;
      END
   END din0[189]
   PIN din0[190]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  681.5425 0.0 681.6825 0.14 ;
      END
   END din0[190]
   PIN din0[191]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  684.4025 0.0 684.5425 0.14 ;
      END
   END din0[191]
   PIN din0[192]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  687.2625 0.0 687.4025 0.14 ;
      END
   END din0[192]
   PIN din0[193]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  690.1225 0.0 690.2625 0.14 ;
      END
   END din0[193]
   PIN din0[194]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  692.9825 0.0 693.1225 0.14 ;
      END
   END din0[194]
   PIN din0[195]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  695.8425 0.0 695.9825 0.14 ;
      END
   END din0[195]
   PIN din0[196]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  698.7025 0.0 698.8425 0.14 ;
      END
   END din0[196]
   PIN din0[197]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  701.5625 0.0 701.7025 0.14 ;
      END
   END din0[197]
   PIN din0[198]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  704.4225 0.0 704.5625 0.14 ;
      END
   END din0[198]
   PIN din0[199]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  707.2825 0.0 707.4225 0.14 ;
      END
   END din0[199]
   PIN din0[200]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  710.1425 0.0 710.2825 0.14 ;
      END
   END din0[200]
   PIN din0[201]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  713.0025 0.0 713.1425 0.14 ;
      END
   END din0[201]
   PIN din0[202]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  715.8625 0.0 716.0025 0.14 ;
      END
   END din0[202]
   PIN din0[203]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  718.7225 0.0 718.8625 0.14 ;
      END
   END din0[203]
   PIN din0[204]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  721.5825 0.0 721.7225 0.14 ;
      END
   END din0[204]
   PIN din0[205]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  724.4425 0.0 724.5825 0.14 ;
      END
   END din0[205]
   PIN din0[206]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  727.3025 0.0 727.4425 0.14 ;
      END
   END din0[206]
   PIN din0[207]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  730.1625 0.0 730.3025 0.14 ;
      END
   END din0[207]
   PIN din0[208]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  733.0225 0.0 733.1625 0.14 ;
      END
   END din0[208]
   PIN din0[209]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  735.8825 0.0 736.0225 0.14 ;
      END
   END din0[209]
   PIN din0[210]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  738.7425 0.0 738.8825 0.14 ;
      END
   END din0[210]
   PIN din0[211]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  741.6025 0.0 741.7425 0.14 ;
      END
   END din0[211]
   PIN din0[212]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  744.4625 0.0 744.6025 0.14 ;
      END
   END din0[212]
   PIN din0[213]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  747.3225 0.0 747.4625 0.14 ;
      END
   END din0[213]
   PIN din0[214]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  750.1825 0.0 750.3225 0.14 ;
      END
   END din0[214]
   PIN din0[215]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  753.0425 0.0 753.1825 0.14 ;
      END
   END din0[215]
   PIN din0[216]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  755.9025 0.0 756.0425 0.14 ;
      END
   END din0[216]
   PIN din0[217]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  758.7625 0.0 758.9025 0.14 ;
      END
   END din0[217]
   PIN din0[218]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  761.6225 0.0 761.7625 0.14 ;
      END
   END din0[218]
   PIN din0[219]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  764.4825 0.0 764.6225 0.14 ;
      END
   END din0[219]
   PIN din0[220]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  767.3425 0.0 767.4825 0.14 ;
      END
   END din0[220]
   PIN din0[221]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  770.2025 0.0 770.3425 0.14 ;
      END
   END din0[221]
   PIN din0[222]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  773.0625 0.0 773.2025 0.14 ;
      END
   END din0[222]
   PIN din0[223]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  775.9225 0.0 776.0625 0.14 ;
      END
   END din0[223]
   PIN din0[224]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  778.7825 0.0 778.9225 0.14 ;
      END
   END din0[224]
   PIN din0[225]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  781.6425 0.0 781.7825 0.14 ;
      END
   END din0[225]
   PIN din0[226]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  784.5025 0.0 784.6425 0.14 ;
      END
   END din0[226]
   PIN din0[227]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  787.3625 0.0 787.5025 0.14 ;
      END
   END din0[227]
   PIN din0[228]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  790.2225 0.0 790.3625 0.14 ;
      END
   END din0[228]
   PIN din0[229]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  793.0825 0.0 793.2225 0.14 ;
      END
   END din0[229]
   PIN din0[230]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  795.9425 0.0 796.0825 0.14 ;
      END
   END din0[230]
   PIN din0[231]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  798.8025 0.0 798.9425 0.14 ;
      END
   END din0[231]
   PIN din0[232]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  801.6625 0.0 801.8025 0.14 ;
      END
   END din0[232]
   PIN din0[233]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  804.5225 0.0 804.6625 0.14 ;
      END
   END din0[233]
   PIN din0[234]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  807.3825 0.0 807.5225 0.14 ;
      END
   END din0[234]
   PIN din0[235]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  810.2425 0.0 810.3825 0.14 ;
      END
   END din0[235]
   PIN din0[236]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  813.1025 0.0 813.2425 0.14 ;
      END
   END din0[236]
   PIN din0[237]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  815.9625 0.0 816.1025 0.14 ;
      END
   END din0[237]
   PIN din0[238]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  818.8225 0.0 818.9625 0.14 ;
      END
   END din0[238]
   PIN din0[239]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  821.6825 0.0 821.8225 0.14 ;
      END
   END din0[239]
   PIN din0[240]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  824.5425 0.0 824.6825 0.14 ;
      END
   END din0[240]
   PIN din0[241]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  827.4025 0.0 827.5425 0.14 ;
      END
   END din0[241]
   PIN din0[242]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  830.2625 0.0 830.4025 0.14 ;
      END
   END din0[242]
   PIN din0[243]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  833.1225 0.0 833.2625 0.14 ;
      END
   END din0[243]
   PIN din0[244]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  835.9825 0.0 836.1225 0.14 ;
      END
   END din0[244]
   PIN din0[245]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  838.8425 0.0 838.9825 0.14 ;
      END
   END din0[245]
   PIN din0[246]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  841.7025 0.0 841.8425 0.14 ;
      END
   END din0[246]
   PIN din0[247]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  844.5625 0.0 844.7025 0.14 ;
      END
   END din0[247]
   PIN din0[248]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  847.4225 0.0 847.5625 0.14 ;
      END
   END din0[248]
   PIN din0[249]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  850.2825 0.0 850.4225 0.14 ;
      END
   END din0[249]
   PIN din0[250]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  853.1425 0.0 853.2825 0.14 ;
      END
   END din0[250]
   PIN din0[251]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  856.0025 0.0 856.1425 0.14 ;
      END
   END din0[251]
   PIN din0[252]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  858.8625 0.0 859.0025 0.14 ;
      END
   END din0[252]
   PIN din0[253]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  861.7225 0.0 861.8625 0.14 ;
      END
   END din0[253]
   PIN din0[254]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  864.5825 0.0 864.7225 0.14 ;
      END
   END din0[254]
   PIN din0[255]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  867.4425 0.0 867.5825 0.14 ;
      END
   END din0[255]
   PIN din0[256]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  870.3025 0.0 870.4425 0.14 ;
      END
   END din0[256]
   PIN din0[257]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  873.1625 0.0 873.3025 0.14 ;
      END
   END din0[257]
   PIN din0[258]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  876.0225 0.0 876.1625 0.14 ;
      END
   END din0[258]
   PIN din0[259]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  878.8825 0.0 879.0225 0.14 ;
      END
   END din0[259]
   PIN din0[260]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  881.7425 0.0 881.8825 0.14 ;
      END
   END din0[260]
   PIN din0[261]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  884.6025 0.0 884.7425 0.14 ;
      END
   END din0[261]
   PIN din0[262]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  887.4625 0.0 887.6025 0.14 ;
      END
   END din0[262]
   PIN din0[263]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  890.3225 0.0 890.4625 0.14 ;
      END
   END din0[263]
   PIN din0[264]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  893.1825 0.0 893.3225 0.14 ;
      END
   END din0[264]
   PIN din0[265]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  896.0425 0.0 896.1825 0.14 ;
      END
   END din0[265]
   PIN din0[266]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  898.9025 0.0 899.0425 0.14 ;
      END
   END din0[266]
   PIN din0[267]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  901.7625 0.0 901.9025 0.14 ;
      END
   END din0[267]
   PIN din0[268]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  904.6225 0.0 904.7625 0.14 ;
      END
   END din0[268]
   PIN din0[269]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  907.4825 0.0 907.6225 0.14 ;
      END
   END din0[269]
   PIN din0[270]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  910.3425 0.0 910.4825 0.14 ;
      END
   END din0[270]
   PIN din0[271]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  913.2025 0.0 913.3425 0.14 ;
      END
   END din0[271]
   PIN din0[272]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  916.0625 0.0 916.2025 0.14 ;
      END
   END din0[272]
   PIN din0[273]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  918.9225 0.0 919.0625 0.14 ;
      END
   END din0[273]
   PIN din0[274]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  921.7825 0.0 921.9225 0.14 ;
      END
   END din0[274]
   PIN din0[275]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  924.6425 0.0 924.7825 0.14 ;
      END
   END din0[275]
   PIN din0[276]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  927.5025 0.0 927.6425 0.14 ;
      END
   END din0[276]
   PIN din0[277]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  930.3625 0.0 930.5025 0.14 ;
      END
   END din0[277]
   PIN din0[278]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  933.2225 0.0 933.3625 0.14 ;
      END
   END din0[278]
   PIN din0[279]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  936.0825 0.0 936.2225 0.14 ;
      END
   END din0[279]
   PIN din0[280]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  938.9425 0.0 939.0825 0.14 ;
      END
   END din0[280]
   PIN din0[281]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  941.8025 0.0 941.9425 0.14 ;
      END
   END din0[281]
   PIN din0[282]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  944.6625 0.0 944.8025 0.14 ;
      END
   END din0[282]
   PIN din0[283]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  947.5225 0.0 947.6625 0.14 ;
      END
   END din0[283]
   PIN din0[284]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  950.3825 0.0 950.5225 0.14 ;
      END
   END din0[284]
   PIN din0[285]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  953.2425 0.0 953.3825 0.14 ;
      END
   END din0[285]
   PIN din0[286]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  956.1025 0.0 956.2425 0.14 ;
      END
   END din0[286]
   PIN din0[287]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  958.9625 0.0 959.1025 0.14 ;
      END
   END din0[287]
   PIN din0[288]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  961.8225 0.0 961.9625 0.14 ;
      END
   END din0[288]
   PIN din0[289]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  964.6825 0.0 964.8225 0.14 ;
      END
   END din0[289]
   PIN din0[290]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  967.5425 0.0 967.6825 0.14 ;
      END
   END din0[290]
   PIN din0[291]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  970.4025 0.0 970.5425 0.14 ;
      END
   END din0[291]
   PIN din0[292]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  973.2625 0.0 973.4025 0.14 ;
      END
   END din0[292]
   PIN din0[293]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  976.1225 0.0 976.2625 0.14 ;
      END
   END din0[293]
   PIN din0[294]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  978.9825 0.0 979.1225 0.14 ;
      END
   END din0[294]
   PIN din0[295]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  981.8425 0.0 981.9825 0.14 ;
      END
   END din0[295]
   PIN din0[296]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  984.7025 0.0 984.8425 0.14 ;
      END
   END din0[296]
   PIN din0[297]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  987.5625 0.0 987.7025 0.14 ;
      END
   END din0[297]
   PIN din0[298]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  990.4225 0.0 990.5625 0.14 ;
      END
   END din0[298]
   PIN din0[299]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  993.2825 0.0 993.4225 0.14 ;
      END
   END din0[299]
   PIN din0[300]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  996.1425 0.0 996.2825 0.14 ;
      END
   END din0[300]
   PIN din0[301]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  999.0025 0.0 999.1425 0.14 ;
      END
   END din0[301]
   PIN din0[302]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1001.8625 0.0 1002.0025 0.14 ;
      END
   END din0[302]
   PIN din0[303]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1004.7225 0.0 1004.8625 0.14 ;
      END
   END din0[303]
   PIN din0[304]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1007.5825 0.0 1007.7225 0.14 ;
      END
   END din0[304]
   PIN din0[305]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1010.4425 0.0 1010.5825 0.14 ;
      END
   END din0[305]
   PIN din0[306]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1013.3025 0.0 1013.4425 0.14 ;
      END
   END din0[306]
   PIN din0[307]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1016.1625 0.0 1016.3025 0.14 ;
      END
   END din0[307]
   PIN din0[308]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1019.0225 0.0 1019.1625 0.14 ;
      END
   END din0[308]
   PIN din0[309]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1021.8825 0.0 1022.0225 0.14 ;
      END
   END din0[309]
   PIN din0[310]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1024.7425 0.0 1024.8825 0.14 ;
      END
   END din0[310]
   PIN din0[311]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1027.6025 0.0 1027.7425 0.14 ;
      END
   END din0[311]
   PIN din0[312]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1030.4625 0.0 1030.6025 0.14 ;
      END
   END din0[312]
   PIN din0[313]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1033.3225 0.0 1033.4625 0.14 ;
      END
   END din0[313]
   PIN din0[314]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1036.1825 0.0 1036.3225 0.14 ;
      END
   END din0[314]
   PIN din0[315]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1039.0425 0.0 1039.1825 0.14 ;
      END
   END din0[315]
   PIN din0[316]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1041.9025 0.0 1042.0425 0.14 ;
      END
   END din0[316]
   PIN din0[317]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1044.7625 0.0 1044.9025 0.14 ;
      END
   END din0[317]
   PIN din0[318]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1047.6225 0.0 1047.7625 0.14 ;
      END
   END din0[318]
   PIN din0[319]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1050.4825 0.0 1050.6225 0.14 ;
      END
   END din0[319]
   PIN din0[320]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1053.3425 0.0 1053.4825 0.14 ;
      END
   END din0[320]
   PIN din0[321]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1056.2025 0.0 1056.3425 0.14 ;
      END
   END din0[321]
   PIN din0[322]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1059.0625 0.0 1059.2025 0.14 ;
      END
   END din0[322]
   PIN din0[323]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1061.9225 0.0 1062.0625 0.14 ;
      END
   END din0[323]
   PIN din0[324]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1064.7825 0.0 1064.9225 0.14 ;
      END
   END din0[324]
   PIN din0[325]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1067.6425 0.0 1067.7825 0.14 ;
      END
   END din0[325]
   PIN din0[326]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1070.5025 0.0 1070.6425 0.14 ;
      END
   END din0[326]
   PIN din0[327]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1073.3625 0.0 1073.5025 0.14 ;
      END
   END din0[327]
   PIN din0[328]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1076.2225 0.0 1076.3625 0.14 ;
      END
   END din0[328]
   PIN din0[329]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1079.0825 0.0 1079.2225 0.14 ;
      END
   END din0[329]
   PIN din0[330]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1081.9425 0.0 1082.0825 0.14 ;
      END
   END din0[330]
   PIN din0[331]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1084.8025 0.0 1084.9425 0.14 ;
      END
   END din0[331]
   PIN din0[332]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1087.6625 0.0 1087.8025 0.14 ;
      END
   END din0[332]
   PIN din0[333]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1090.5225 0.0 1090.6625 0.14 ;
      END
   END din0[333]
   PIN din0[334]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1093.3825 0.0 1093.5225 0.14 ;
      END
   END din0[334]
   PIN din0[335]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1096.2425 0.0 1096.3825 0.14 ;
      END
   END din0[335]
   PIN din0[336]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1099.1025 0.0 1099.2425 0.14 ;
      END
   END din0[336]
   PIN din0[337]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1101.9625 0.0 1102.1025 0.14 ;
      END
   END din0[337]
   PIN din0[338]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1104.8225 0.0 1104.9625 0.14 ;
      END
   END din0[338]
   PIN din0[339]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1107.6825 0.0 1107.8225 0.14 ;
      END
   END din0[339]
   PIN din0[340]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1110.5425 0.0 1110.6825 0.14 ;
      END
   END din0[340]
   PIN din0[341]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1113.4025 0.0 1113.5425 0.14 ;
      END
   END din0[341]
   PIN din0[342]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1116.2625 0.0 1116.4025 0.14 ;
      END
   END din0[342]
   PIN din0[343]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1119.1225 0.0 1119.2625 0.14 ;
      END
   END din0[343]
   PIN din0[344]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1121.9825 0.0 1122.1225 0.14 ;
      END
   END din0[344]
   PIN din0[345]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1124.8425 0.0 1124.9825 0.14 ;
      END
   END din0[345]
   PIN din0[346]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1127.7025 0.0 1127.8425 0.14 ;
      END
   END din0[346]
   PIN din0[347]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1130.5625 0.0 1130.7025 0.14 ;
      END
   END din0[347]
   PIN din0[348]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1133.4225 0.0 1133.5625 0.14 ;
      END
   END din0[348]
   PIN din0[349]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1136.2825 0.0 1136.4225 0.14 ;
      END
   END din0[349]
   PIN din0[350]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1139.1425 0.0 1139.2825 0.14 ;
      END
   END din0[350]
   PIN din0[351]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1142.0025 0.0 1142.1425 0.14 ;
      END
   END din0[351]
   PIN din0[352]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1144.8625 0.0 1145.0025 0.14 ;
      END
   END din0[352]
   PIN din0[353]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1147.7225 0.0 1147.8625 0.14 ;
      END
   END din0[353]
   PIN din0[354]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1150.5825 0.0 1150.7225 0.14 ;
      END
   END din0[354]
   PIN din0[355]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1153.4425 0.0 1153.5825 0.14 ;
      END
   END din0[355]
   PIN din0[356]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1156.3025 0.0 1156.4425 0.14 ;
      END
   END din0[356]
   PIN din0[357]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1159.1625 0.0 1159.3025 0.14 ;
      END
   END din0[357]
   PIN din0[358]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1162.0225 0.0 1162.1625 0.14 ;
      END
   END din0[358]
   PIN din0[359]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1164.8825 0.0 1165.0225 0.14 ;
      END
   END din0[359]
   PIN din0[360]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1167.7425 0.0 1167.8825 0.14 ;
      END
   END din0[360]
   PIN din0[361]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1170.6025 0.0 1170.7425 0.14 ;
      END
   END din0[361]
   PIN din0[362]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1173.4625 0.0 1173.6025 0.14 ;
      END
   END din0[362]
   PIN din0[363]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1176.3225 0.0 1176.4625 0.14 ;
      END
   END din0[363]
   PIN din0[364]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1179.1825 0.0 1179.3225 0.14 ;
      END
   END din0[364]
   PIN din0[365]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1182.0425 0.0 1182.1825 0.14 ;
      END
   END din0[365]
   PIN din0[366]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1184.9025 0.0 1185.0425 0.14 ;
      END
   END din0[366]
   PIN din0[367]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1187.7625 0.0 1187.9025 0.14 ;
      END
   END din0[367]
   PIN din0[368]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1190.6225 0.0 1190.7625 0.14 ;
      END
   END din0[368]
   PIN din0[369]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1193.4825 0.0 1193.6225 0.14 ;
      END
   END din0[369]
   PIN din0[370]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1196.3425 0.0 1196.4825 0.14 ;
      END
   END din0[370]
   PIN din0[371]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1199.2025 0.0 1199.3425 0.14 ;
      END
   END din0[371]
   PIN din0[372]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1202.0625 0.0 1202.2025 0.14 ;
      END
   END din0[372]
   PIN din0[373]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1204.9225 0.0 1205.0625 0.14 ;
      END
   END din0[373]
   PIN din0[374]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1207.7825 0.0 1207.9225 0.14 ;
      END
   END din0[374]
   PIN din0[375]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1210.6425 0.0 1210.7825 0.14 ;
      END
   END din0[375]
   PIN din0[376]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1213.5025 0.0 1213.6425 0.14 ;
      END
   END din0[376]
   PIN din0[377]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1216.3625 0.0 1216.5025 0.14 ;
      END
   END din0[377]
   PIN din0[378]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1219.2225 0.0 1219.3625 0.14 ;
      END
   END din0[378]
   PIN din0[379]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1222.0825 0.0 1222.2225 0.14 ;
      END
   END din0[379]
   PIN din0[380]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1224.9425 0.0 1225.0825 0.14 ;
      END
   END din0[380]
   PIN din0[381]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1227.8025 0.0 1227.9425 0.14 ;
      END
   END din0[381]
   PIN din0[382]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1230.6625 0.0 1230.8025 0.14 ;
      END
   END din0[382]
   PIN din0[383]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1233.5225 0.0 1233.6625 0.14 ;
      END
   END din0[383]
   PIN din0[384]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1236.3825 0.0 1236.5225 0.14 ;
      END
   END din0[384]
   PIN din0[385]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1239.2425 0.0 1239.3825 0.14 ;
      END
   END din0[385]
   PIN din0[386]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1242.1025 0.0 1242.2425 0.14 ;
      END
   END din0[386]
   PIN din0[387]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1244.9625 0.0 1245.1025 0.14 ;
      END
   END din0[387]
   PIN din0[388]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1247.8225 0.0 1247.9625 0.14 ;
      END
   END din0[388]
   PIN din0[389]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1250.6825 0.0 1250.8225 0.14 ;
      END
   END din0[389]
   PIN din0[390]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1253.5425 0.0 1253.6825 0.14 ;
      END
   END din0[390]
   PIN din0[391]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1256.4025 0.0 1256.5425 0.14 ;
      END
   END din0[391]
   PIN din0[392]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1259.2625 0.0 1259.4025 0.14 ;
      END
   END din0[392]
   PIN din0[393]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1262.1225 0.0 1262.2625 0.14 ;
      END
   END din0[393]
   PIN din0[394]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1264.9825 0.0 1265.1225 0.14 ;
      END
   END din0[394]
   PIN din0[395]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1267.8425 0.0 1267.9825 0.14 ;
      END
   END din0[395]
   PIN din0[396]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1270.7025 0.0 1270.8425 0.14 ;
      END
   END din0[396]
   PIN din0[397]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1273.5625 0.0 1273.7025 0.14 ;
      END
   END din0[397]
   PIN din0[398]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1276.4225 0.0 1276.5625 0.14 ;
      END
   END din0[398]
   PIN din0[399]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1279.2825 0.0 1279.4225 0.14 ;
      END
   END din0[399]
   PIN din0[400]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1282.1425 0.0 1282.2825 0.14 ;
      END
   END din0[400]
   PIN din0[401]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1285.0025 0.0 1285.1425 0.14 ;
      END
   END din0[401]
   PIN din0[402]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1287.8625 0.0 1288.0025 0.14 ;
      END
   END din0[402]
   PIN din0[403]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1290.7225 0.0 1290.8625 0.14 ;
      END
   END din0[403]
   PIN din0[404]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1293.5825 0.0 1293.7225 0.14 ;
      END
   END din0[404]
   PIN din0[405]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1296.4425 0.0 1296.5825 0.14 ;
      END
   END din0[405]
   PIN din0[406]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1299.3025 0.0 1299.4425 0.14 ;
      END
   END din0[406]
   PIN din0[407]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1302.1625 0.0 1302.3025 0.14 ;
      END
   END din0[407]
   PIN din0[408]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1305.0225 0.0 1305.1625 0.14 ;
      END
   END din0[408]
   PIN din0[409]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1307.8825 0.0 1308.0225 0.14 ;
      END
   END din0[409]
   PIN din0[410]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1310.7425 0.0 1310.8825 0.14 ;
      END
   END din0[410]
   PIN din0[411]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1313.6025 0.0 1313.7425 0.14 ;
      END
   END din0[411]
   PIN din0[412]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1316.4625 0.0 1316.6025 0.14 ;
      END
   END din0[412]
   PIN din0[413]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1319.3225 0.0 1319.4625 0.14 ;
      END
   END din0[413]
   PIN din0[414]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1322.1825 0.0 1322.3225 0.14 ;
      END
   END din0[414]
   PIN din0[415]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1325.0425 0.0 1325.1825 0.14 ;
      END
   END din0[415]
   PIN din0[416]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1327.9025 0.0 1328.0425 0.14 ;
      END
   END din0[416]
   PIN din0[417]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1330.7625 0.0 1330.9025 0.14 ;
      END
   END din0[417]
   PIN din0[418]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1333.6225 0.0 1333.7625 0.14 ;
      END
   END din0[418]
   PIN din0[419]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1336.4825 0.0 1336.6225 0.14 ;
      END
   END din0[419]
   PIN din0[420]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1339.3425 0.0 1339.4825 0.14 ;
      END
   END din0[420]
   PIN din0[421]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1342.2025 0.0 1342.3425 0.14 ;
      END
   END din0[421]
   PIN din0[422]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1345.0625 0.0 1345.2025 0.14 ;
      END
   END din0[422]
   PIN din0[423]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1347.9225 0.0 1348.0625 0.14 ;
      END
   END din0[423]
   PIN din0[424]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1350.7825 0.0 1350.9225 0.14 ;
      END
   END din0[424]
   PIN din0[425]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1353.6425 0.0 1353.7825 0.14 ;
      END
   END din0[425]
   PIN din0[426]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1356.5025 0.0 1356.6425 0.14 ;
      END
   END din0[426]
   PIN din0[427]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1359.3625 0.0 1359.5025 0.14 ;
      END
   END din0[427]
   PIN din0[428]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1362.2225 0.0 1362.3625 0.14 ;
      END
   END din0[428]
   PIN din0[429]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1365.0825 0.0 1365.2225 0.14 ;
      END
   END din0[429]
   PIN din0[430]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1367.9425 0.0 1368.0825 0.14 ;
      END
   END din0[430]
   PIN din0[431]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1370.8025 0.0 1370.9425 0.14 ;
      END
   END din0[431]
   PIN din0[432]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1373.6625 0.0 1373.8025 0.14 ;
      END
   END din0[432]
   PIN din0[433]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1376.5225 0.0 1376.6625 0.14 ;
      END
   END din0[433]
   PIN din0[434]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1379.3825 0.0 1379.5225 0.14 ;
      END
   END din0[434]
   PIN din0[435]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1382.2425 0.0 1382.3825 0.14 ;
      END
   END din0[435]
   PIN din0[436]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1385.1025 0.0 1385.2425 0.14 ;
      END
   END din0[436]
   PIN din0[437]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1387.9625 0.0 1388.1025 0.14 ;
      END
   END din0[437]
   PIN din0[438]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1390.8225 0.0 1390.9625 0.14 ;
      END
   END din0[438]
   PIN din0[439]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1393.6825 0.0 1393.8225 0.14 ;
      END
   END din0[439]
   PIN din0[440]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1396.5425 0.0 1396.6825 0.14 ;
      END
   END din0[440]
   PIN din0[441]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1399.4025 0.0 1399.5425 0.14 ;
      END
   END din0[441]
   PIN din0[442]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1402.2625 0.0 1402.4025 0.14 ;
      END
   END din0[442]
   PIN din0[443]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1405.1225 0.0 1405.2625 0.14 ;
      END
   END din0[443]
   PIN din0[444]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1407.9825 0.0 1408.1225 0.14 ;
      END
   END din0[444]
   PIN din0[445]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1410.8425 0.0 1410.9825 0.14 ;
      END
   END din0[445]
   PIN din0[446]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1413.7025 0.0 1413.8425 0.14 ;
      END
   END din0[446]
   PIN din0[447]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1416.5625 0.0 1416.7025 0.14 ;
      END
   END din0[447]
   PIN din0[448]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1419.4225 0.0 1419.5625 0.14 ;
      END
   END din0[448]
   PIN din0[449]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1422.2825 0.0 1422.4225 0.14 ;
      END
   END din0[449]
   PIN din0[450]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1425.1425 0.0 1425.2825 0.14 ;
      END
   END din0[450]
   PIN din0[451]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1428.0025 0.0 1428.1425 0.14 ;
      END
   END din0[451]
   PIN din0[452]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1430.8625 0.0 1431.0025 0.14 ;
      END
   END din0[452]
   PIN din0[453]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1433.7225 0.0 1433.8625 0.14 ;
      END
   END din0[453]
   PIN din0[454]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1436.5825 0.0 1436.7225 0.14 ;
      END
   END din0[454]
   PIN din0[455]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1439.4425 0.0 1439.5825 0.14 ;
      END
   END din0[455]
   PIN din0[456]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1442.3025 0.0 1442.4425 0.14 ;
      END
   END din0[456]
   PIN din0[457]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1445.1625 0.0 1445.3025 0.14 ;
      END
   END din0[457]
   PIN din0[458]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1448.0225 0.0 1448.1625 0.14 ;
      END
   END din0[458]
   PIN din0[459]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1450.8825 0.0 1451.0225 0.14 ;
      END
   END din0[459]
   PIN din0[460]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1453.7425 0.0 1453.8825 0.14 ;
      END
   END din0[460]
   PIN din0[461]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1456.6025 0.0 1456.7425 0.14 ;
      END
   END din0[461]
   PIN din0[462]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1459.4625 0.0 1459.6025 0.14 ;
      END
   END din0[462]
   PIN din0[463]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1462.3225 0.0 1462.4625 0.14 ;
      END
   END din0[463]
   PIN din0[464]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1465.1825 0.0 1465.3225 0.14 ;
      END
   END din0[464]
   PIN din0[465]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1468.0425 0.0 1468.1825 0.14 ;
      END
   END din0[465]
   PIN din0[466]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1470.9025 0.0 1471.0425 0.14 ;
      END
   END din0[466]
   PIN din0[467]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1473.7625 0.0 1473.9025 0.14 ;
      END
   END din0[467]
   PIN din0[468]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1476.6225 0.0 1476.7625 0.14 ;
      END
   END din0[468]
   PIN din0[469]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1479.4825 0.0 1479.6225 0.14 ;
      END
   END din0[469]
   PIN din0[470]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1482.3425 0.0 1482.4825 0.14 ;
      END
   END din0[470]
   PIN din0[471]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1485.2025 0.0 1485.3425 0.14 ;
      END
   END din0[471]
   PIN din0[472]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1488.0625 0.0 1488.2025 0.14 ;
      END
   END din0[472]
   PIN din0[473]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1490.9225 0.0 1491.0625 0.14 ;
      END
   END din0[473]
   PIN din0[474]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1493.7825 0.0 1493.9225 0.14 ;
      END
   END din0[474]
   PIN din0[475]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1496.6425 0.0 1496.7825 0.14 ;
      END
   END din0[475]
   PIN din0[476]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1499.5025 0.0 1499.6425 0.14 ;
      END
   END din0[476]
   PIN din0[477]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1502.3625 0.0 1502.5025 0.14 ;
      END
   END din0[477]
   PIN din0[478]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1505.2225 0.0 1505.3625 0.14 ;
      END
   END din0[478]
   PIN din0[479]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1508.0825 0.0 1508.2225 0.14 ;
      END
   END din0[479]
   PIN din0[480]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1510.9425 0.0 1511.0825 0.14 ;
      END
   END din0[480]
   PIN din0[481]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1513.8025 0.0 1513.9425 0.14 ;
      END
   END din0[481]
   PIN din0[482]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1516.6625 0.0 1516.8025 0.14 ;
      END
   END din0[482]
   PIN din0[483]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1519.5225 0.0 1519.6625 0.14 ;
      END
   END din0[483]
   PIN din0[484]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1522.3825 0.0 1522.5225 0.14 ;
      END
   END din0[484]
   PIN din0[485]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1525.2425 0.0 1525.3825 0.14 ;
      END
   END din0[485]
   PIN din0[486]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1528.1025 0.0 1528.2425 0.14 ;
      END
   END din0[486]
   PIN din0[487]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1530.9625 0.0 1531.1025 0.14 ;
      END
   END din0[487]
   PIN din0[488]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1533.8225 0.0 1533.9625 0.14 ;
      END
   END din0[488]
   PIN din0[489]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1536.6825 0.0 1536.8225 0.14 ;
      END
   END din0[489]
   PIN din0[490]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1539.5425 0.0 1539.6825 0.14 ;
      END
   END din0[490]
   PIN din0[491]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1542.4025 0.0 1542.5425 0.14 ;
      END
   END din0[491]
   PIN din0[492]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1545.2625 0.0 1545.4025 0.14 ;
      END
   END din0[492]
   PIN din0[493]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1548.1225 0.0 1548.2625 0.14 ;
      END
   END din0[493]
   PIN din0[494]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1550.9825 0.0 1551.1225 0.14 ;
      END
   END din0[494]
   PIN din0[495]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1553.8425 0.0 1553.9825 0.14 ;
      END
   END din0[495]
   PIN din0[496]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1556.7025 0.0 1556.8425 0.14 ;
      END
   END din0[496]
   PIN din0[497]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1559.5625 0.0 1559.7025 0.14 ;
      END
   END din0[497]
   PIN din0[498]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1562.4225 0.0 1562.5625 0.14 ;
      END
   END din0[498]
   PIN din0[499]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1565.2825 0.0 1565.4225 0.14 ;
      END
   END din0[499]
   PIN din0[500]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1568.1425 0.0 1568.2825 0.14 ;
      END
   END din0[500]
   PIN din0[501]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1571.0025 0.0 1571.1425 0.14 ;
      END
   END din0[501]
   PIN din0[502]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1573.8625 0.0 1574.0025 0.14 ;
      END
   END din0[502]
   PIN din0[503]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1576.7225 0.0 1576.8625 0.14 ;
      END
   END din0[503]
   PIN din0[504]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1579.5825 0.0 1579.7225 0.14 ;
      END
   END din0[504]
   PIN din0[505]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1582.4425 0.0 1582.5825 0.14 ;
      END
   END din0[505]
   PIN din0[506]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1585.3025 0.0 1585.4425 0.14 ;
      END
   END din0[506]
   PIN din0[507]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1588.1625 0.0 1588.3025 0.14 ;
      END
   END din0[507]
   PIN din0[508]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1591.0225 0.0 1591.1625 0.14 ;
      END
   END din0[508]
   PIN din0[509]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1593.8825 0.0 1594.0225 0.14 ;
      END
   END din0[509]
   PIN din0[510]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1596.7425 0.0 1596.8825 0.14 ;
      END
   END din0[510]
   PIN din0[511]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1599.6025 0.0 1599.7425 0.14 ;
      END
   END din0[511]
   PIN din0[512]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1602.4625 0.0 1602.6025 0.14 ;
      END
   END din0[512]
   PIN din0[513]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1605.3225 0.0 1605.4625 0.14 ;
      END
   END din0[513]
   PIN din0[514]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1608.1825 0.0 1608.3225 0.14 ;
      END
   END din0[514]
   PIN din0[515]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1611.0425 0.0 1611.1825 0.14 ;
      END
   END din0[515]
   PIN din0[516]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1613.9025 0.0 1614.0425 0.14 ;
      END
   END din0[516]
   PIN din0[517]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1616.7625 0.0 1616.9025 0.14 ;
      END
   END din0[517]
   PIN din0[518]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1619.6225 0.0 1619.7625 0.14 ;
      END
   END din0[518]
   PIN din0[519]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1622.4825 0.0 1622.6225 0.14 ;
      END
   END din0[519]
   PIN din0[520]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1625.3425 0.0 1625.4825 0.14 ;
      END
   END din0[520]
   PIN din0[521]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1628.2025 0.0 1628.3425 0.14 ;
      END
   END din0[521]
   PIN din0[522]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1631.0625 0.0 1631.2025 0.14 ;
      END
   END din0[522]
   PIN din0[523]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1633.9225 0.0 1634.0625 0.14 ;
      END
   END din0[523]
   PIN din0[524]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1636.7825 0.0 1636.9225 0.14 ;
      END
   END din0[524]
   PIN din0[525]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1639.6425 0.0 1639.7825 0.14 ;
      END
   END din0[525]
   PIN din0[526]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1642.5025 0.0 1642.6425 0.14 ;
      END
   END din0[526]
   PIN din0[527]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1645.3625 0.0 1645.5025 0.14 ;
      END
   END din0[527]
   PIN din0[528]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1648.2225 0.0 1648.3625 0.14 ;
      END
   END din0[528]
   PIN din0[529]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1651.0825 0.0 1651.2225 0.14 ;
      END
   END din0[529]
   PIN din0[530]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1653.9425 0.0 1654.0825 0.14 ;
      END
   END din0[530]
   PIN din0[531]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1656.8025 0.0 1656.9425 0.14 ;
      END
   END din0[531]
   PIN din0[532]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1659.6625 0.0 1659.8025 0.14 ;
      END
   END din0[532]
   PIN din0[533]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1662.5225 0.0 1662.6625 0.14 ;
      END
   END din0[533]
   PIN din0[534]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1665.3825 0.0 1665.5225 0.14 ;
      END
   END din0[534]
   PIN din0[535]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1668.2425 0.0 1668.3825 0.14 ;
      END
   END din0[535]
   PIN din0[536]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1671.1025 0.0 1671.2425 0.14 ;
      END
   END din0[536]
   PIN din0[537]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1673.9625 0.0 1674.1025 0.14 ;
      END
   END din0[537]
   PIN din0[538]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1676.8225 0.0 1676.9625 0.14 ;
      END
   END din0[538]
   PIN din0[539]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1679.6825 0.0 1679.8225 0.14 ;
      END
   END din0[539]
   PIN din0[540]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1682.5425 0.0 1682.6825 0.14 ;
      END
   END din0[540]
   PIN din0[541]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1685.4025 0.0 1685.5425 0.14 ;
      END
   END din0[541]
   PIN din0[542]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1688.2625 0.0 1688.4025 0.14 ;
      END
   END din0[542]
   PIN din0[543]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1691.1225 0.0 1691.2625 0.14 ;
      END
   END din0[543]
   PIN din0[544]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1693.9825 0.0 1694.1225 0.14 ;
      END
   END din0[544]
   PIN din0[545]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1696.8425 0.0 1696.9825 0.14 ;
      END
   END din0[545]
   PIN din0[546]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1699.7025 0.0 1699.8425 0.14 ;
      END
   END din0[546]
   PIN din0[547]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1702.5625 0.0 1702.7025 0.14 ;
      END
   END din0[547]
   PIN din0[548]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1705.4225 0.0 1705.5625 0.14 ;
      END
   END din0[548]
   PIN din0[549]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1708.2825 0.0 1708.4225 0.14 ;
      END
   END din0[549]
   PIN din0[550]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1711.1425 0.0 1711.2825 0.14 ;
      END
   END din0[550]
   PIN din0[551]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1714.0025 0.0 1714.1425 0.14 ;
      END
   END din0[551]
   PIN din0[552]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1716.8625 0.0 1717.0025 0.14 ;
      END
   END din0[552]
   PIN din0[553]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1719.7225 0.0 1719.8625 0.14 ;
      END
   END din0[553]
   PIN din0[554]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1722.5825 0.0 1722.7225 0.14 ;
      END
   END din0[554]
   PIN din0[555]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1725.4425 0.0 1725.5825 0.14 ;
      END
   END din0[555]
   PIN din0[556]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1728.3025 0.0 1728.4425 0.14 ;
      END
   END din0[556]
   PIN din0[557]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1731.1625 0.0 1731.3025 0.14 ;
      END
   END din0[557]
   PIN din0[558]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1734.0225 0.0 1734.1625 0.14 ;
      END
   END din0[558]
   PIN din0[559]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1736.8825 0.0 1737.0225 0.14 ;
      END
   END din0[559]
   PIN din0[560]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1739.7425 0.0 1739.8825 0.14 ;
      END
   END din0[560]
   PIN din0[561]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1742.6025 0.0 1742.7425 0.14 ;
      END
   END din0[561]
   PIN din0[562]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1745.4625 0.0 1745.6025 0.14 ;
      END
   END din0[562]
   PIN din0[563]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1748.3225 0.0 1748.4625 0.14 ;
      END
   END din0[563]
   PIN din0[564]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1751.1825 0.0 1751.3225 0.14 ;
      END
   END din0[564]
   PIN din0[565]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1754.0425 0.0 1754.1825 0.14 ;
      END
   END din0[565]
   PIN din0[566]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1756.9025 0.0 1757.0425 0.14 ;
      END
   END din0[566]
   PIN din0[567]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1759.7625 0.0 1759.9025 0.14 ;
      END
   END din0[567]
   PIN din0[568]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1762.6225 0.0 1762.7625 0.14 ;
      END
   END din0[568]
   PIN din0[569]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1765.4825 0.0 1765.6225 0.14 ;
      END
   END din0[569]
   PIN din0[570]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1768.3425 0.0 1768.4825 0.14 ;
      END
   END din0[570]
   PIN din0[571]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1771.2025 0.0 1771.3425 0.14 ;
      END
   END din0[571]
   PIN din0[572]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1774.0625 0.0 1774.2025 0.14 ;
      END
   END din0[572]
   PIN din0[573]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1776.9225 0.0 1777.0625 0.14 ;
      END
   END din0[573]
   PIN din0[574]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1779.7825 0.0 1779.9225 0.14 ;
      END
   END din0[574]
   PIN din0[575]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1782.6425 0.0 1782.7825 0.14 ;
      END
   END din0[575]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  132.995 192.83 133.135 192.97 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  131.855 192.83 131.995 192.97 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  132.71 192.83 132.85 192.97 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  132.425 192.83 132.565 192.97 ;
      END
   END addr0[3]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  891.63 192.83 891.77 192.97 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  891.345 192.83 891.485 192.97 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  892.2 192.83 892.34 192.97 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  891.63 192.83 891.77 192.97 ;
      END
   END addr1[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 88.18 0.14 88.32 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1020.6925 192.83 1020.8325 192.97 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 88.415 0.14 88.555 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  1014.495 192.83 1014.635 192.97 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  173.5575 192.83 173.6975 192.97 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  174.7325 192.83 174.8725 192.97 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  175.9075 192.83 176.0475 192.97 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  177.0825 192.83 177.2225 192.97 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  178.2575 192.83 178.3975 192.97 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  179.4325 192.83 179.5725 192.97 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  180.6075 192.83 180.7475 192.97 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  181.7825 192.83 181.9225 192.97 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  182.9575 192.83 183.0975 192.97 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  184.1325 192.83 184.2725 192.97 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  185.3075 192.83 185.4475 192.97 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  186.4825 192.83 186.6225 192.97 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  187.6575 192.83 187.7975 192.97 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  188.8325 192.83 188.9725 192.97 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  190.0075 192.83 190.1475 192.97 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  191.1825 192.83 191.3225 192.97 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  192.3575 192.83 192.4975 192.97 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  193.5325 192.83 193.6725 192.97 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  194.7075 192.83 194.8475 192.97 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  195.8825 192.83 196.0225 192.97 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  197.0575 192.83 197.1975 192.97 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  198.2325 192.83 198.3725 192.97 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  199.4075 192.83 199.5475 192.97 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  200.5825 192.83 200.7225 192.97 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  201.7575 192.83 201.8975 192.97 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  202.9325 192.83 203.0725 192.97 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  204.1075 192.83 204.2475 192.97 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  205.2825 192.83 205.4225 192.97 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  206.4575 192.83 206.5975 192.97 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  207.6325 192.83 207.7725 192.97 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  208.8075 192.83 208.9475 192.97 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  209.9825 192.83 210.1225 192.97 ;
      END
   END dout1[31]
   PIN dout1[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  211.1575 192.83 211.2975 192.97 ;
      END
   END dout1[32]
   PIN dout1[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  212.3325 192.83 212.4725 192.97 ;
      END
   END dout1[33]
   PIN dout1[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  213.5075 192.83 213.6475 192.97 ;
      END
   END dout1[34]
   PIN dout1[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  214.6825 192.83 214.8225 192.97 ;
      END
   END dout1[35]
   PIN dout1[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  215.8575 192.83 215.9975 192.97 ;
      END
   END dout1[36]
   PIN dout1[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  217.0325 192.83 217.1725 192.97 ;
      END
   END dout1[37]
   PIN dout1[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  218.2075 192.83 218.3475 192.97 ;
      END
   END dout1[38]
   PIN dout1[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  219.3825 192.83 219.5225 192.97 ;
      END
   END dout1[39]
   PIN dout1[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  220.5575 192.83 220.6975 192.97 ;
      END
   END dout1[40]
   PIN dout1[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  221.7325 192.83 221.8725 192.97 ;
      END
   END dout1[41]
   PIN dout1[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  222.9075 192.83 223.0475 192.97 ;
      END
   END dout1[42]
   PIN dout1[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  224.0825 192.83 224.2225 192.97 ;
      END
   END dout1[43]
   PIN dout1[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  225.2575 192.83 225.3975 192.97 ;
      END
   END dout1[44]
   PIN dout1[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  226.4325 192.83 226.5725 192.97 ;
      END
   END dout1[45]
   PIN dout1[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  227.6075 192.83 227.7475 192.97 ;
      END
   END dout1[46]
   PIN dout1[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  228.7825 192.83 228.9225 192.97 ;
      END
   END dout1[47]
   PIN dout1[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  229.9575 192.83 230.0975 192.97 ;
      END
   END dout1[48]
   PIN dout1[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  231.1325 192.83 231.2725 192.97 ;
      END
   END dout1[49]
   PIN dout1[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  232.3075 192.83 232.4475 192.97 ;
      END
   END dout1[50]
   PIN dout1[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  233.4825 192.83 233.6225 192.97 ;
      END
   END dout1[51]
   PIN dout1[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  234.6575 192.83 234.7975 192.97 ;
      END
   END dout1[52]
   PIN dout1[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  235.8325 192.83 235.9725 192.97 ;
      END
   END dout1[53]
   PIN dout1[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  237.0075 192.83 237.1475 192.97 ;
      END
   END dout1[54]
   PIN dout1[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  238.1825 192.83 238.3225 192.97 ;
      END
   END dout1[55]
   PIN dout1[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  239.3575 192.83 239.4975 192.97 ;
      END
   END dout1[56]
   PIN dout1[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  240.5325 192.83 240.6725 192.97 ;
      END
   END dout1[57]
   PIN dout1[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  241.7075 192.83 241.8475 192.97 ;
      END
   END dout1[58]
   PIN dout1[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  242.8825 192.83 243.0225 192.97 ;
      END
   END dout1[59]
   PIN dout1[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  244.0575 192.83 244.1975 192.97 ;
      END
   END dout1[60]
   PIN dout1[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  245.2325 192.83 245.3725 192.97 ;
      END
   END dout1[61]
   PIN dout1[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  246.4075 192.83 246.5475 192.97 ;
      END
   END dout1[62]
   PIN dout1[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  247.5825 192.83 247.7225 192.97 ;
      END
   END dout1[63]
   PIN dout1[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  248.7575 192.83 248.8975 192.97 ;
      END
   END dout1[64]
   PIN dout1[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  249.9325 192.83 250.0725 192.97 ;
      END
   END dout1[65]
   PIN dout1[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  251.1075 192.83 251.2475 192.97 ;
      END
   END dout1[66]
   PIN dout1[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  252.2825 192.83 252.4225 192.97 ;
      END
   END dout1[67]
   PIN dout1[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  253.4575 192.83 253.5975 192.97 ;
      END
   END dout1[68]
   PIN dout1[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  254.6325 192.83 254.7725 192.97 ;
      END
   END dout1[69]
   PIN dout1[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  255.8075 192.83 255.9475 192.97 ;
      END
   END dout1[70]
   PIN dout1[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  256.9825 192.83 257.1225 192.97 ;
      END
   END dout1[71]
   PIN dout1[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  258.1575 192.83 258.2975 192.97 ;
      END
   END dout1[72]
   PIN dout1[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  259.3325 192.83 259.4725 192.97 ;
      END
   END dout1[73]
   PIN dout1[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  260.5075 192.83 260.6475 192.97 ;
      END
   END dout1[74]
   PIN dout1[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  261.6825 192.83 261.8225 192.97 ;
      END
   END dout1[75]
   PIN dout1[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  262.8575 192.83 262.9975 192.97 ;
      END
   END dout1[76]
   PIN dout1[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  264.0325 192.83 264.1725 192.97 ;
      END
   END dout1[77]
   PIN dout1[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  265.2075 192.83 265.3475 192.97 ;
      END
   END dout1[78]
   PIN dout1[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  266.3825 192.83 266.5225 192.97 ;
      END
   END dout1[79]
   PIN dout1[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  267.5575 192.83 267.6975 192.97 ;
      END
   END dout1[80]
   PIN dout1[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  268.7325 192.83 268.8725 192.97 ;
      END
   END dout1[81]
   PIN dout1[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  269.9075 192.83 270.0475 192.97 ;
      END
   END dout1[82]
   PIN dout1[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  271.0825 192.83 271.2225 192.97 ;
      END
   END dout1[83]
   PIN dout1[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  272.2575 192.83 272.3975 192.97 ;
      END
   END dout1[84]
   PIN dout1[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  273.4325 192.83 273.5725 192.97 ;
      END
   END dout1[85]
   PIN dout1[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  274.6075 192.83 274.7475 192.97 ;
      END
   END dout1[86]
   PIN dout1[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  275.7825 192.83 275.9225 192.97 ;
      END
   END dout1[87]
   PIN dout1[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  276.9575 192.83 277.0975 192.97 ;
      END
   END dout1[88]
   PIN dout1[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  278.1325 192.83 278.2725 192.97 ;
      END
   END dout1[89]
   PIN dout1[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  279.3075 192.83 279.4475 192.97 ;
      END
   END dout1[90]
   PIN dout1[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  280.4825 192.83 280.6225 192.97 ;
      END
   END dout1[91]
   PIN dout1[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  281.6575 192.83 281.7975 192.97 ;
      END
   END dout1[92]
   PIN dout1[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  282.8325 192.83 282.9725 192.97 ;
      END
   END dout1[93]
   PIN dout1[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  284.0075 192.83 284.1475 192.97 ;
      END
   END dout1[94]
   PIN dout1[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  285.1825 192.83 285.3225 192.97 ;
      END
   END dout1[95]
   PIN dout1[96]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  286.3575 192.83 286.4975 192.97 ;
      END
   END dout1[96]
   PIN dout1[97]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  287.5325 192.83 287.6725 192.97 ;
      END
   END dout1[97]
   PIN dout1[98]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  288.7075 192.83 288.8475 192.97 ;
      END
   END dout1[98]
   PIN dout1[99]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  289.8825 192.83 290.0225 192.97 ;
      END
   END dout1[99]
   PIN dout1[100]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  291.0575 192.83 291.1975 192.97 ;
      END
   END dout1[100]
   PIN dout1[101]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  292.2325 192.83 292.3725 192.97 ;
      END
   END dout1[101]
   PIN dout1[102]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  293.4075 192.83 293.5475 192.97 ;
      END
   END dout1[102]
   PIN dout1[103]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  294.5825 192.83 294.7225 192.97 ;
      END
   END dout1[103]
   PIN dout1[104]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  295.7575 192.83 295.8975 192.97 ;
      END
   END dout1[104]
   PIN dout1[105]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  296.9325 192.83 297.0725 192.97 ;
      END
   END dout1[105]
   PIN dout1[106]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  298.1075 192.83 298.2475 192.97 ;
      END
   END dout1[106]
   PIN dout1[107]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  299.2825 192.83 299.4225 192.97 ;
      END
   END dout1[107]
   PIN dout1[108]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  300.4575 192.83 300.5975 192.97 ;
      END
   END dout1[108]
   PIN dout1[109]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  301.6325 192.83 301.7725 192.97 ;
      END
   END dout1[109]
   PIN dout1[110]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  302.8075 192.83 302.9475 192.97 ;
      END
   END dout1[110]
   PIN dout1[111]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  303.9825 192.83 304.1225 192.97 ;
      END
   END dout1[111]
   PIN dout1[112]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  305.1575 192.83 305.2975 192.97 ;
      END
   END dout1[112]
   PIN dout1[113]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  306.3325 192.83 306.4725 192.97 ;
      END
   END dout1[113]
   PIN dout1[114]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  307.5075 192.83 307.6475 192.97 ;
      END
   END dout1[114]
   PIN dout1[115]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  308.6825 192.83 308.8225 192.97 ;
      END
   END dout1[115]
   PIN dout1[116]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  309.8575 192.83 309.9975 192.97 ;
      END
   END dout1[116]
   PIN dout1[117]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  311.0325 192.83 311.1725 192.97 ;
      END
   END dout1[117]
   PIN dout1[118]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  312.2075 192.83 312.3475 192.97 ;
      END
   END dout1[118]
   PIN dout1[119]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  313.3825 192.83 313.5225 192.97 ;
      END
   END dout1[119]
   PIN dout1[120]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  314.5575 192.83 314.6975 192.97 ;
      END
   END dout1[120]
   PIN dout1[121]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  315.7325 192.83 315.8725 192.97 ;
      END
   END dout1[121]
   PIN dout1[122]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  316.9075 192.83 317.0475 192.97 ;
      END
   END dout1[122]
   PIN dout1[123]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  318.0825 192.83 318.2225 192.97 ;
      END
   END dout1[123]
   PIN dout1[124]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  319.2575 192.83 319.3975 192.97 ;
      END
   END dout1[124]
   PIN dout1[125]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  320.4325 192.83 320.5725 192.97 ;
      END
   END dout1[125]
   PIN dout1[126]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  321.6075 192.83 321.7475 192.97 ;
      END
   END dout1[126]
   PIN dout1[127]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  322.7825 192.83 322.9225 192.97 ;
      END
   END dout1[127]
   PIN dout1[128]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  323.9575 192.83 324.0975 192.97 ;
      END
   END dout1[128]
   PIN dout1[129]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  325.1325 192.83 325.2725 192.97 ;
      END
   END dout1[129]
   PIN dout1[130]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  326.3075 192.83 326.4475 192.97 ;
      END
   END dout1[130]
   PIN dout1[131]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  327.4825 192.83 327.6225 192.97 ;
      END
   END dout1[131]
   PIN dout1[132]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  328.6575 192.83 328.7975 192.97 ;
      END
   END dout1[132]
   PIN dout1[133]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  329.8325 192.83 329.9725 192.97 ;
      END
   END dout1[133]
   PIN dout1[134]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  331.0075 192.83 331.1475 192.97 ;
      END
   END dout1[134]
   PIN dout1[135]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  332.1825 192.83 332.3225 192.97 ;
      END
   END dout1[135]
   PIN dout1[136]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  333.3575 192.83 333.4975 192.97 ;
      END
   END dout1[136]
   PIN dout1[137]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  334.5325 192.83 334.6725 192.97 ;
      END
   END dout1[137]
   PIN dout1[138]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  335.7075 192.83 335.8475 192.97 ;
      END
   END dout1[138]
   PIN dout1[139]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  336.8825 192.83 337.0225 192.97 ;
      END
   END dout1[139]
   PIN dout1[140]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  338.0575 192.83 338.1975 192.97 ;
      END
   END dout1[140]
   PIN dout1[141]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  339.2325 192.83 339.3725 192.97 ;
      END
   END dout1[141]
   PIN dout1[142]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  340.4075 192.83 340.5475 192.97 ;
      END
   END dout1[142]
   PIN dout1[143]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  341.5825 192.83 341.7225 192.97 ;
      END
   END dout1[143]
   PIN dout1[144]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  342.7575 192.83 342.8975 192.97 ;
      END
   END dout1[144]
   PIN dout1[145]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  343.9325 192.83 344.0725 192.97 ;
      END
   END dout1[145]
   PIN dout1[146]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  345.1075 192.83 345.2475 192.97 ;
      END
   END dout1[146]
   PIN dout1[147]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  346.2825 192.83 346.4225 192.97 ;
      END
   END dout1[147]
   PIN dout1[148]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  347.4575 192.83 347.5975 192.97 ;
      END
   END dout1[148]
   PIN dout1[149]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  348.6325 192.83 348.7725 192.97 ;
      END
   END dout1[149]
   PIN dout1[150]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  349.8075 192.83 349.9475 192.97 ;
      END
   END dout1[150]
   PIN dout1[151]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  350.9825 192.83 351.1225 192.97 ;
      END
   END dout1[151]
   PIN dout1[152]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  352.1575 192.83 352.2975 192.97 ;
      END
   END dout1[152]
   PIN dout1[153]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  353.3325 192.83 353.4725 192.97 ;
      END
   END dout1[153]
   PIN dout1[154]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  354.5075 192.83 354.6475 192.97 ;
      END
   END dout1[154]
   PIN dout1[155]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  355.6825 192.83 355.8225 192.97 ;
      END
   END dout1[155]
   PIN dout1[156]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  356.8575 192.83 356.9975 192.97 ;
      END
   END dout1[156]
   PIN dout1[157]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  358.0325 192.83 358.1725 192.97 ;
      END
   END dout1[157]
   PIN dout1[158]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  359.2075 192.83 359.3475 192.97 ;
      END
   END dout1[158]
   PIN dout1[159]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  360.3825 192.83 360.5225 192.97 ;
      END
   END dout1[159]
   PIN dout1[160]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  361.5575 192.83 361.6975 192.97 ;
      END
   END dout1[160]
   PIN dout1[161]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  362.7325 192.83 362.8725 192.97 ;
      END
   END dout1[161]
   PIN dout1[162]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  363.9075 192.83 364.0475 192.97 ;
      END
   END dout1[162]
   PIN dout1[163]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  365.0825 192.83 365.2225 192.97 ;
      END
   END dout1[163]
   PIN dout1[164]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  366.2575 192.83 366.3975 192.97 ;
      END
   END dout1[164]
   PIN dout1[165]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  367.4325 192.83 367.5725 192.97 ;
      END
   END dout1[165]
   PIN dout1[166]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  368.6075 192.83 368.7475 192.97 ;
      END
   END dout1[166]
   PIN dout1[167]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  369.7825 192.83 369.9225 192.97 ;
      END
   END dout1[167]
   PIN dout1[168]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  370.9575 192.83 371.0975 192.97 ;
      END
   END dout1[168]
   PIN dout1[169]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  372.1325 192.83 372.2725 192.97 ;
      END
   END dout1[169]
   PIN dout1[170]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  373.3075 192.83 373.4475 192.97 ;
      END
   END dout1[170]
   PIN dout1[171]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  374.4825 192.83 374.6225 192.97 ;
      END
   END dout1[171]
   PIN dout1[172]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  375.6575 192.83 375.7975 192.97 ;
      END
   END dout1[172]
   PIN dout1[173]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  376.8325 192.83 376.9725 192.97 ;
      END
   END dout1[173]
   PIN dout1[174]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  378.0075 192.83 378.1475 192.97 ;
      END
   END dout1[174]
   PIN dout1[175]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  379.1825 192.83 379.3225 192.97 ;
      END
   END dout1[175]
   PIN dout1[176]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  380.3575 192.83 380.4975 192.97 ;
      END
   END dout1[176]
   PIN dout1[177]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  381.5325 192.83 381.6725 192.97 ;
      END
   END dout1[177]
   PIN dout1[178]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  382.7075 192.83 382.8475 192.97 ;
      END
   END dout1[178]
   PIN dout1[179]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  383.8825 192.83 384.0225 192.97 ;
      END
   END dout1[179]
   PIN dout1[180]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  385.0575 192.83 385.1975 192.97 ;
      END
   END dout1[180]
   PIN dout1[181]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  386.2325 192.83 386.3725 192.97 ;
      END
   END dout1[181]
   PIN dout1[182]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  387.4075 192.83 387.5475 192.97 ;
      END
   END dout1[182]
   PIN dout1[183]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  388.5825 192.83 388.7225 192.97 ;
      END
   END dout1[183]
   PIN dout1[184]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  389.7575 192.83 389.8975 192.97 ;
      END
   END dout1[184]
   PIN dout1[185]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  390.9325 192.83 391.0725 192.97 ;
      END
   END dout1[185]
   PIN dout1[186]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  392.1075 192.83 392.2475 192.97 ;
      END
   END dout1[186]
   PIN dout1[187]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  393.2825 192.83 393.4225 192.97 ;
      END
   END dout1[187]
   PIN dout1[188]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  394.4575 192.83 394.5975 192.97 ;
      END
   END dout1[188]
   PIN dout1[189]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  395.6325 192.83 395.7725 192.97 ;
      END
   END dout1[189]
   PIN dout1[190]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  396.8075 192.83 396.9475 192.97 ;
      END
   END dout1[190]
   PIN dout1[191]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  397.9825 192.83 398.1225 192.97 ;
      END
   END dout1[191]
   PIN dout1[192]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  399.1575 192.83 399.2975 192.97 ;
      END
   END dout1[192]
   PIN dout1[193]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  400.3325 192.83 400.4725 192.97 ;
      END
   END dout1[193]
   PIN dout1[194]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  401.5075 192.83 401.6475 192.97 ;
      END
   END dout1[194]
   PIN dout1[195]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  402.6825 192.83 402.8225 192.97 ;
      END
   END dout1[195]
   PIN dout1[196]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  403.8575 192.83 403.9975 192.97 ;
      END
   END dout1[196]
   PIN dout1[197]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  405.0325 192.83 405.1725 192.97 ;
      END
   END dout1[197]
   PIN dout1[198]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  406.2075 192.83 406.3475 192.97 ;
      END
   END dout1[198]
   PIN dout1[199]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  407.3825 192.83 407.5225 192.97 ;
      END
   END dout1[199]
   PIN dout1[200]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  408.5575 192.83 408.6975 192.97 ;
      END
   END dout1[200]
   PIN dout1[201]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  409.7325 192.83 409.8725 192.97 ;
      END
   END dout1[201]
   PIN dout1[202]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  410.9075 192.83 411.0475 192.97 ;
      END
   END dout1[202]
   PIN dout1[203]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  412.0825 192.83 412.2225 192.97 ;
      END
   END dout1[203]
   PIN dout1[204]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  413.2575 192.83 413.3975 192.97 ;
      END
   END dout1[204]
   PIN dout1[205]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  414.4325 192.83 414.5725 192.97 ;
      END
   END dout1[205]
   PIN dout1[206]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  415.6075 192.83 415.7475 192.97 ;
      END
   END dout1[206]
   PIN dout1[207]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  416.7825 192.83 416.9225 192.97 ;
      END
   END dout1[207]
   PIN dout1[208]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  417.9575 192.83 418.0975 192.97 ;
      END
   END dout1[208]
   PIN dout1[209]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  419.1325 192.83 419.2725 192.97 ;
      END
   END dout1[209]
   PIN dout1[210]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  420.3075 192.83 420.4475 192.97 ;
      END
   END dout1[210]
   PIN dout1[211]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  421.4825 192.83 421.6225 192.97 ;
      END
   END dout1[211]
   PIN dout1[212]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  422.6575 192.83 422.7975 192.97 ;
      END
   END dout1[212]
   PIN dout1[213]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  423.8325 192.83 423.9725 192.97 ;
      END
   END dout1[213]
   PIN dout1[214]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  425.0075 192.83 425.1475 192.97 ;
      END
   END dout1[214]
   PIN dout1[215]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  426.1825 192.83 426.3225 192.97 ;
      END
   END dout1[215]
   PIN dout1[216]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  427.3575 192.83 427.4975 192.97 ;
      END
   END dout1[216]
   PIN dout1[217]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  428.5325 192.83 428.6725 192.97 ;
      END
   END dout1[217]
   PIN dout1[218]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  429.7075 192.83 429.8475 192.97 ;
      END
   END dout1[218]
   PIN dout1[219]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  430.8825 192.83 431.0225 192.97 ;
      END
   END dout1[219]
   PIN dout1[220]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  432.0575 192.83 432.1975 192.97 ;
      END
   END dout1[220]
   PIN dout1[221]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  433.2325 192.83 433.3725 192.97 ;
      END
   END dout1[221]
   PIN dout1[222]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  434.4075 192.83 434.5475 192.97 ;
      END
   END dout1[222]
   PIN dout1[223]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  435.5825 192.83 435.7225 192.97 ;
      END
   END dout1[223]
   PIN dout1[224]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  436.7575 192.83 436.8975 192.97 ;
      END
   END dout1[224]
   PIN dout1[225]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  437.9325 192.83 438.0725 192.97 ;
      END
   END dout1[225]
   PIN dout1[226]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  439.1075 192.83 439.2475 192.97 ;
      END
   END dout1[226]
   PIN dout1[227]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  440.2825 192.83 440.4225 192.97 ;
      END
   END dout1[227]
   PIN dout1[228]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  441.4575 192.83 441.5975 192.97 ;
      END
   END dout1[228]
   PIN dout1[229]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  442.6325 192.83 442.7725 192.97 ;
      END
   END dout1[229]
   PIN dout1[230]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  443.8075 192.83 443.9475 192.97 ;
      END
   END dout1[230]
   PIN dout1[231]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  444.9825 192.83 445.1225 192.97 ;
      END
   END dout1[231]
   PIN dout1[232]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  446.1575 192.83 446.2975 192.97 ;
      END
   END dout1[232]
   PIN dout1[233]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  447.3325 192.83 447.4725 192.97 ;
      END
   END dout1[233]
   PIN dout1[234]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  448.5075 192.83 448.6475 192.97 ;
      END
   END dout1[234]
   PIN dout1[235]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  449.6825 192.83 449.8225 192.97 ;
      END
   END dout1[235]
   PIN dout1[236]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  450.8575 192.83 450.9975 192.97 ;
      END
   END dout1[236]
   PIN dout1[237]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  452.0325 192.83 452.1725 192.97 ;
      END
   END dout1[237]
   PIN dout1[238]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  453.2075 192.83 453.3475 192.97 ;
      END
   END dout1[238]
   PIN dout1[239]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  454.3825 192.83 454.5225 192.97 ;
      END
   END dout1[239]
   PIN dout1[240]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  455.5575 192.83 455.6975 192.97 ;
      END
   END dout1[240]
   PIN dout1[241]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  456.7325 192.83 456.8725 192.97 ;
      END
   END dout1[241]
   PIN dout1[242]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  457.9075 192.83 458.0475 192.97 ;
      END
   END dout1[242]
   PIN dout1[243]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  459.0825 192.83 459.2225 192.97 ;
      END
   END dout1[243]
   PIN dout1[244]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  460.2575 192.83 460.3975 192.97 ;
      END
   END dout1[244]
   PIN dout1[245]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  461.4325 192.83 461.5725 192.97 ;
      END
   END dout1[245]
   PIN dout1[246]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  462.6075 192.83 462.7475 192.97 ;
      END
   END dout1[246]
   PIN dout1[247]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  463.7825 192.83 463.9225 192.97 ;
      END
   END dout1[247]
   PIN dout1[248]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  464.9575 192.83 465.0975 192.97 ;
      END
   END dout1[248]
   PIN dout1[249]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  466.1325 192.83 466.2725 192.97 ;
      END
   END dout1[249]
   PIN dout1[250]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  467.3075 192.83 467.4475 192.97 ;
      END
   END dout1[250]
   PIN dout1[251]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  468.4825 192.83 468.6225 192.97 ;
      END
   END dout1[251]
   PIN dout1[252]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  469.6575 192.83 469.7975 192.97 ;
      END
   END dout1[252]
   PIN dout1[253]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  470.8325 192.83 470.9725 192.97 ;
      END
   END dout1[253]
   PIN dout1[254]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  472.0075 192.83 472.1475 192.97 ;
      END
   END dout1[254]
   PIN dout1[255]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  473.1825 192.83 473.3225 192.97 ;
      END
   END dout1[255]
   PIN dout1[256]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  474.3575 192.83 474.4975 192.97 ;
      END
   END dout1[256]
   PIN dout1[257]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  475.5325 192.83 475.6725 192.97 ;
      END
   END dout1[257]
   PIN dout1[258]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  476.7075 192.83 476.8475 192.97 ;
      END
   END dout1[258]
   PIN dout1[259]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  477.8825 192.83 478.0225 192.97 ;
      END
   END dout1[259]
   PIN dout1[260]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  479.0575 192.83 479.1975 192.97 ;
      END
   END dout1[260]
   PIN dout1[261]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  480.2325 192.83 480.3725 192.97 ;
      END
   END dout1[261]
   PIN dout1[262]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  481.4075 192.83 481.5475 192.97 ;
      END
   END dout1[262]
   PIN dout1[263]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  482.5825 192.83 482.7225 192.97 ;
      END
   END dout1[263]
   PIN dout1[264]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  483.7575 192.83 483.8975 192.97 ;
      END
   END dout1[264]
   PIN dout1[265]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  484.9325 192.83 485.0725 192.97 ;
      END
   END dout1[265]
   PIN dout1[266]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  486.1075 192.83 486.2475 192.97 ;
      END
   END dout1[266]
   PIN dout1[267]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  487.2825 192.83 487.4225 192.97 ;
      END
   END dout1[267]
   PIN dout1[268]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  488.4575 192.83 488.5975 192.97 ;
      END
   END dout1[268]
   PIN dout1[269]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  489.6325 192.83 489.7725 192.97 ;
      END
   END dout1[269]
   PIN dout1[270]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  490.8075 192.83 490.9475 192.97 ;
      END
   END dout1[270]
   PIN dout1[271]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  491.9825 192.83 492.1225 192.97 ;
      END
   END dout1[271]
   PIN dout1[272]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  493.1575 192.83 493.2975 192.97 ;
      END
   END dout1[272]
   PIN dout1[273]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  494.3325 192.83 494.4725 192.97 ;
      END
   END dout1[273]
   PIN dout1[274]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  495.5075 192.83 495.6475 192.97 ;
      END
   END dout1[274]
   PIN dout1[275]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  496.6825 192.83 496.8225 192.97 ;
      END
   END dout1[275]
   PIN dout1[276]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  497.8575 192.83 497.9975 192.97 ;
      END
   END dout1[276]
   PIN dout1[277]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  499.0325 192.83 499.1725 192.97 ;
      END
   END dout1[277]
   PIN dout1[278]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  500.2075 192.83 500.3475 192.97 ;
      END
   END dout1[278]
   PIN dout1[279]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  501.3825 192.83 501.5225 192.97 ;
      END
   END dout1[279]
   PIN dout1[280]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  502.5575 192.83 502.6975 192.97 ;
      END
   END dout1[280]
   PIN dout1[281]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  503.7325 192.83 503.8725 192.97 ;
      END
   END dout1[281]
   PIN dout1[282]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  504.9075 192.83 505.0475 192.97 ;
      END
   END dout1[282]
   PIN dout1[283]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  506.0825 192.83 506.2225 192.97 ;
      END
   END dout1[283]
   PIN dout1[284]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  507.2575 192.83 507.3975 192.97 ;
      END
   END dout1[284]
   PIN dout1[285]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  508.4325 192.83 508.5725 192.97 ;
      END
   END dout1[285]
   PIN dout1[286]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  509.6075 192.83 509.7475 192.97 ;
      END
   END dout1[286]
   PIN dout1[287]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  510.7825 192.83 510.9225 192.97 ;
      END
   END dout1[287]
   PIN dout1[288]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  511.9575 192.83 512.0975 192.97 ;
      END
   END dout1[288]
   PIN dout1[289]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  513.1325 192.83 513.2725 192.97 ;
      END
   END dout1[289]
   PIN dout1[290]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  514.3075 192.83 514.4475 192.97 ;
      END
   END dout1[290]
   PIN dout1[291]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  515.4825 192.83 515.6225 192.97 ;
      END
   END dout1[291]
   PIN dout1[292]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  516.6575 192.83 516.7975 192.97 ;
      END
   END dout1[292]
   PIN dout1[293]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  517.8325 192.83 517.9725 192.97 ;
      END
   END dout1[293]
   PIN dout1[294]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  519.0075 192.83 519.1475 192.97 ;
      END
   END dout1[294]
   PIN dout1[295]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  520.1825 192.83 520.3225 192.97 ;
      END
   END dout1[295]
   PIN dout1[296]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  521.3575 192.83 521.4975 192.97 ;
      END
   END dout1[296]
   PIN dout1[297]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  522.5325 192.83 522.6725 192.97 ;
      END
   END dout1[297]
   PIN dout1[298]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  523.7075 192.83 523.8475 192.97 ;
      END
   END dout1[298]
   PIN dout1[299]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  524.8825 192.83 525.0225 192.97 ;
      END
   END dout1[299]
   PIN dout1[300]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  526.0575 192.83 526.1975 192.97 ;
      END
   END dout1[300]
   PIN dout1[301]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  527.2325 192.83 527.3725 192.97 ;
      END
   END dout1[301]
   PIN dout1[302]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  528.4075 192.83 528.5475 192.97 ;
      END
   END dout1[302]
   PIN dout1[303]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  529.5825 192.83 529.7225 192.97 ;
      END
   END dout1[303]
   PIN dout1[304]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  530.7575 192.83 530.8975 192.97 ;
      END
   END dout1[304]
   PIN dout1[305]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  531.9325 192.83 532.0725 192.97 ;
      END
   END dout1[305]
   PIN dout1[306]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  533.1075 192.83 533.2475 192.97 ;
      END
   END dout1[306]
   PIN dout1[307]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  534.2825 192.83 534.4225 192.97 ;
      END
   END dout1[307]
   PIN dout1[308]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  535.4575 192.83 535.5975 192.97 ;
      END
   END dout1[308]
   PIN dout1[309]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  536.6325 192.83 536.7725 192.97 ;
      END
   END dout1[309]
   PIN dout1[310]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  537.8075 192.83 537.9475 192.97 ;
      END
   END dout1[310]
   PIN dout1[311]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  538.9825 192.83 539.1225 192.97 ;
      END
   END dout1[311]
   PIN dout1[312]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  540.1575 192.83 540.2975 192.97 ;
      END
   END dout1[312]
   PIN dout1[313]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  541.3325 192.83 541.4725 192.97 ;
      END
   END dout1[313]
   PIN dout1[314]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  542.5075 192.83 542.6475 192.97 ;
      END
   END dout1[314]
   PIN dout1[315]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  543.6825 192.83 543.8225 192.97 ;
      END
   END dout1[315]
   PIN dout1[316]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  544.8575 192.83 544.9975 192.97 ;
      END
   END dout1[316]
   PIN dout1[317]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  546.0325 192.83 546.1725 192.97 ;
      END
   END dout1[317]
   PIN dout1[318]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  547.2075 192.83 547.3475 192.97 ;
      END
   END dout1[318]
   PIN dout1[319]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  548.3825 192.83 548.5225 192.97 ;
      END
   END dout1[319]
   PIN dout1[320]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  549.5575 192.83 549.6975 192.97 ;
      END
   END dout1[320]
   PIN dout1[321]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  550.7325 192.83 550.8725 192.97 ;
      END
   END dout1[321]
   PIN dout1[322]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  551.9075 192.83 552.0475 192.97 ;
      END
   END dout1[322]
   PIN dout1[323]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  553.0825 192.83 553.2225 192.97 ;
      END
   END dout1[323]
   PIN dout1[324]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  554.2575 192.83 554.3975 192.97 ;
      END
   END dout1[324]
   PIN dout1[325]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  555.4325 192.83 555.5725 192.97 ;
      END
   END dout1[325]
   PIN dout1[326]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  556.6075 192.83 556.7475 192.97 ;
      END
   END dout1[326]
   PIN dout1[327]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  557.7825 192.83 557.9225 192.97 ;
      END
   END dout1[327]
   PIN dout1[328]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  558.9575 192.83 559.0975 192.97 ;
      END
   END dout1[328]
   PIN dout1[329]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  560.1325 192.83 560.2725 192.97 ;
      END
   END dout1[329]
   PIN dout1[330]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  561.3075 192.83 561.4475 192.97 ;
      END
   END dout1[330]
   PIN dout1[331]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  562.4825 192.83 562.6225 192.97 ;
      END
   END dout1[331]
   PIN dout1[332]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  563.6575 192.83 563.7975 192.97 ;
      END
   END dout1[332]
   PIN dout1[333]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  564.8325 192.83 564.9725 192.97 ;
      END
   END dout1[333]
   PIN dout1[334]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  566.0075 192.83 566.1475 192.97 ;
      END
   END dout1[334]
   PIN dout1[335]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  567.1825 192.83 567.3225 192.97 ;
      END
   END dout1[335]
   PIN dout1[336]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  568.3575 192.83 568.4975 192.97 ;
      END
   END dout1[336]
   PIN dout1[337]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  569.5325 192.83 569.6725 192.97 ;
      END
   END dout1[337]
   PIN dout1[338]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  570.7075 192.83 570.8475 192.97 ;
      END
   END dout1[338]
   PIN dout1[339]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  571.8825 192.83 572.0225 192.97 ;
      END
   END dout1[339]
   PIN dout1[340]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  573.0575 192.83 573.1975 192.97 ;
      END
   END dout1[340]
   PIN dout1[341]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  574.2325 192.83 574.3725 192.97 ;
      END
   END dout1[341]
   PIN dout1[342]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  575.4075 192.83 575.5475 192.97 ;
      END
   END dout1[342]
   PIN dout1[343]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  576.5825 192.83 576.7225 192.97 ;
      END
   END dout1[343]
   PIN dout1[344]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  577.7575 192.83 577.8975 192.97 ;
      END
   END dout1[344]
   PIN dout1[345]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  578.9325 192.83 579.0725 192.97 ;
      END
   END dout1[345]
   PIN dout1[346]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  580.1075 192.83 580.2475 192.97 ;
      END
   END dout1[346]
   PIN dout1[347]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  581.2825 192.83 581.4225 192.97 ;
      END
   END dout1[347]
   PIN dout1[348]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  582.4575 192.83 582.5975 192.97 ;
      END
   END dout1[348]
   PIN dout1[349]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  583.6325 192.83 583.7725 192.97 ;
      END
   END dout1[349]
   PIN dout1[350]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  584.8075 192.83 584.9475 192.97 ;
      END
   END dout1[350]
   PIN dout1[351]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  585.9825 192.83 586.1225 192.97 ;
      END
   END dout1[351]
   PIN dout1[352]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  587.1575 192.83 587.2975 192.97 ;
      END
   END dout1[352]
   PIN dout1[353]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  588.3325 192.83 588.4725 192.97 ;
      END
   END dout1[353]
   PIN dout1[354]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  589.5075 192.83 589.6475 192.97 ;
      END
   END dout1[354]
   PIN dout1[355]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  590.6825 192.83 590.8225 192.97 ;
      END
   END dout1[355]
   PIN dout1[356]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  591.8575 192.83 591.9975 192.97 ;
      END
   END dout1[356]
   PIN dout1[357]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  593.0325 192.83 593.1725 192.97 ;
      END
   END dout1[357]
   PIN dout1[358]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  594.2075 192.83 594.3475 192.97 ;
      END
   END dout1[358]
   PIN dout1[359]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  595.3825 192.83 595.5225 192.97 ;
      END
   END dout1[359]
   PIN dout1[360]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  596.5575 192.83 596.6975 192.97 ;
      END
   END dout1[360]
   PIN dout1[361]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  597.7325 192.83 597.8725 192.97 ;
      END
   END dout1[361]
   PIN dout1[362]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  598.9075 192.83 599.0475 192.97 ;
      END
   END dout1[362]
   PIN dout1[363]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  600.0825 192.83 600.2225 192.97 ;
      END
   END dout1[363]
   PIN dout1[364]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  601.2575 192.83 601.3975 192.97 ;
      END
   END dout1[364]
   PIN dout1[365]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  602.4325 192.83 602.5725 192.97 ;
      END
   END dout1[365]
   PIN dout1[366]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  603.6075 192.83 603.7475 192.97 ;
      END
   END dout1[366]
   PIN dout1[367]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  604.7825 192.83 604.9225 192.97 ;
      END
   END dout1[367]
   PIN dout1[368]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  605.9575 192.83 606.0975 192.97 ;
      END
   END dout1[368]
   PIN dout1[369]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  607.1325 192.83 607.2725 192.97 ;
      END
   END dout1[369]
   PIN dout1[370]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  608.3075 192.83 608.4475 192.97 ;
      END
   END dout1[370]
   PIN dout1[371]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  609.4825 192.83 609.6225 192.97 ;
      END
   END dout1[371]
   PIN dout1[372]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  610.6575 192.83 610.7975 192.97 ;
      END
   END dout1[372]
   PIN dout1[373]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  611.8325 192.83 611.9725 192.97 ;
      END
   END dout1[373]
   PIN dout1[374]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  613.0075 192.83 613.1475 192.97 ;
      END
   END dout1[374]
   PIN dout1[375]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  614.1825 192.83 614.3225 192.97 ;
      END
   END dout1[375]
   PIN dout1[376]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  615.3575 192.83 615.4975 192.97 ;
      END
   END dout1[376]
   PIN dout1[377]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  616.5325 192.83 616.6725 192.97 ;
      END
   END dout1[377]
   PIN dout1[378]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  617.7075 192.83 617.8475 192.97 ;
      END
   END dout1[378]
   PIN dout1[379]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  618.8825 192.83 619.0225 192.97 ;
      END
   END dout1[379]
   PIN dout1[380]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  620.0575 192.83 620.1975 192.97 ;
      END
   END dout1[380]
   PIN dout1[381]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  621.2325 192.83 621.3725 192.97 ;
      END
   END dout1[381]
   PIN dout1[382]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  622.4075 192.83 622.5475 192.97 ;
      END
   END dout1[382]
   PIN dout1[383]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  623.5825 192.83 623.7225 192.97 ;
      END
   END dout1[383]
   PIN dout1[384]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  624.7575 192.83 624.8975 192.97 ;
      END
   END dout1[384]
   PIN dout1[385]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  625.9325 192.83 626.0725 192.97 ;
      END
   END dout1[385]
   PIN dout1[386]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  627.1075 192.83 627.2475 192.97 ;
      END
   END dout1[386]
   PIN dout1[387]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  628.2825 192.83 628.4225 192.97 ;
      END
   END dout1[387]
   PIN dout1[388]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  629.4575 192.83 629.5975 192.97 ;
      END
   END dout1[388]
   PIN dout1[389]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  630.6325 192.83 630.7725 192.97 ;
      END
   END dout1[389]
   PIN dout1[390]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  631.8075 192.83 631.9475 192.97 ;
      END
   END dout1[390]
   PIN dout1[391]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  632.9825 192.83 633.1225 192.97 ;
      END
   END dout1[391]
   PIN dout1[392]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  634.1575 192.83 634.2975 192.97 ;
      END
   END dout1[392]
   PIN dout1[393]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  635.3325 192.83 635.4725 192.97 ;
      END
   END dout1[393]
   PIN dout1[394]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  636.5075 192.83 636.6475 192.97 ;
      END
   END dout1[394]
   PIN dout1[395]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  637.6825 192.83 637.8225 192.97 ;
      END
   END dout1[395]
   PIN dout1[396]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  638.8575 192.83 638.9975 192.97 ;
      END
   END dout1[396]
   PIN dout1[397]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  640.0325 192.83 640.1725 192.97 ;
      END
   END dout1[397]
   PIN dout1[398]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  641.2075 192.83 641.3475 192.97 ;
      END
   END dout1[398]
   PIN dout1[399]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  642.3825 192.83 642.5225 192.97 ;
      END
   END dout1[399]
   PIN dout1[400]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  643.5575 192.83 643.6975 192.97 ;
      END
   END dout1[400]
   PIN dout1[401]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  644.7325 192.83 644.8725 192.97 ;
      END
   END dout1[401]
   PIN dout1[402]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  645.9075 192.83 646.0475 192.97 ;
      END
   END dout1[402]
   PIN dout1[403]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  647.0825 192.83 647.2225 192.97 ;
      END
   END dout1[403]
   PIN dout1[404]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  648.2575 192.83 648.3975 192.97 ;
      END
   END dout1[404]
   PIN dout1[405]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  649.4325 192.83 649.5725 192.97 ;
      END
   END dout1[405]
   PIN dout1[406]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  650.6075 192.83 650.7475 192.97 ;
      END
   END dout1[406]
   PIN dout1[407]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  651.7825 192.83 651.9225 192.97 ;
      END
   END dout1[407]
   PIN dout1[408]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  652.9575 192.83 653.0975 192.97 ;
      END
   END dout1[408]
   PIN dout1[409]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  654.1325 192.83 654.2725 192.97 ;
      END
   END dout1[409]
   PIN dout1[410]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  655.3075 192.83 655.4475 192.97 ;
      END
   END dout1[410]
   PIN dout1[411]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  656.4825 192.83 656.6225 192.97 ;
      END
   END dout1[411]
   PIN dout1[412]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  657.6575 192.83 657.7975 192.97 ;
      END
   END dout1[412]
   PIN dout1[413]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  658.8325 192.83 658.9725 192.97 ;
      END
   END dout1[413]
   PIN dout1[414]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  660.0075 192.83 660.1475 192.97 ;
      END
   END dout1[414]
   PIN dout1[415]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  661.1825 192.83 661.3225 192.97 ;
      END
   END dout1[415]
   PIN dout1[416]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  662.3575 192.83 662.4975 192.97 ;
      END
   END dout1[416]
   PIN dout1[417]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  663.5325 192.83 663.6725 192.97 ;
      END
   END dout1[417]
   PIN dout1[418]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  664.7075 192.83 664.8475 192.97 ;
      END
   END dout1[418]
   PIN dout1[419]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  665.8825 192.83 666.0225 192.97 ;
      END
   END dout1[419]
   PIN dout1[420]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  667.0575 192.83 667.1975 192.97 ;
      END
   END dout1[420]
   PIN dout1[421]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  668.2325 192.83 668.3725 192.97 ;
      END
   END dout1[421]
   PIN dout1[422]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  669.4075 192.83 669.5475 192.97 ;
      END
   END dout1[422]
   PIN dout1[423]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  670.5825 192.83 670.7225 192.97 ;
      END
   END dout1[423]
   PIN dout1[424]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  671.7575 192.83 671.8975 192.97 ;
      END
   END dout1[424]
   PIN dout1[425]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  672.9325 192.83 673.0725 192.97 ;
      END
   END dout1[425]
   PIN dout1[426]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  674.1075 192.83 674.2475 192.97 ;
      END
   END dout1[426]
   PIN dout1[427]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  675.2825 192.83 675.4225 192.97 ;
      END
   END dout1[427]
   PIN dout1[428]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  676.4575 192.83 676.5975 192.97 ;
      END
   END dout1[428]
   PIN dout1[429]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  677.6325 192.83 677.7725 192.97 ;
      END
   END dout1[429]
   PIN dout1[430]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  678.8075 192.83 678.9475 192.97 ;
      END
   END dout1[430]
   PIN dout1[431]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  679.9825 192.83 680.1225 192.97 ;
      END
   END dout1[431]
   PIN dout1[432]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  681.1575 192.83 681.2975 192.97 ;
      END
   END dout1[432]
   PIN dout1[433]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  682.3325 192.83 682.4725 192.97 ;
      END
   END dout1[433]
   PIN dout1[434]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  683.5075 192.83 683.6475 192.97 ;
      END
   END dout1[434]
   PIN dout1[435]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  684.6825 192.83 684.8225 192.97 ;
      END
   END dout1[435]
   PIN dout1[436]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  685.8575 192.83 685.9975 192.97 ;
      END
   END dout1[436]
   PIN dout1[437]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  687.0325 192.83 687.1725 192.97 ;
      END
   END dout1[437]
   PIN dout1[438]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  688.2075 192.83 688.3475 192.97 ;
      END
   END dout1[438]
   PIN dout1[439]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  689.3825 192.83 689.5225 192.97 ;
      END
   END dout1[439]
   PIN dout1[440]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  690.5575 192.83 690.6975 192.97 ;
      END
   END dout1[440]
   PIN dout1[441]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  691.7325 192.83 691.8725 192.97 ;
      END
   END dout1[441]
   PIN dout1[442]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  692.9075 192.83 693.0475 192.97 ;
      END
   END dout1[442]
   PIN dout1[443]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  694.0825 192.83 694.2225 192.97 ;
      END
   END dout1[443]
   PIN dout1[444]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  695.2575 192.83 695.3975 192.97 ;
      END
   END dout1[444]
   PIN dout1[445]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  696.4325 192.83 696.5725 192.97 ;
      END
   END dout1[445]
   PIN dout1[446]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  697.6075 192.83 697.7475 192.97 ;
      END
   END dout1[446]
   PIN dout1[447]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  698.7825 192.83 698.9225 192.97 ;
      END
   END dout1[447]
   PIN dout1[448]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  699.9575 192.83 700.0975 192.97 ;
      END
   END dout1[448]
   PIN dout1[449]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  701.1325 192.83 701.2725 192.97 ;
      END
   END dout1[449]
   PIN dout1[450]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  702.3075 192.83 702.4475 192.97 ;
      END
   END dout1[450]
   PIN dout1[451]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  703.4825 192.83 703.6225 192.97 ;
      END
   END dout1[451]
   PIN dout1[452]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  704.6575 192.83 704.7975 192.97 ;
      END
   END dout1[452]
   PIN dout1[453]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  705.8325 192.83 705.9725 192.97 ;
      END
   END dout1[453]
   PIN dout1[454]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  707.0075 192.83 707.1475 192.97 ;
      END
   END dout1[454]
   PIN dout1[455]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  708.1825 192.83 708.3225 192.97 ;
      END
   END dout1[455]
   PIN dout1[456]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  709.3575 192.83 709.4975 192.97 ;
      END
   END dout1[456]
   PIN dout1[457]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  710.5325 192.83 710.6725 192.97 ;
      END
   END dout1[457]
   PIN dout1[458]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  711.7075 192.83 711.8475 192.97 ;
      END
   END dout1[458]
   PIN dout1[459]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  712.8825 192.83 713.0225 192.97 ;
      END
   END dout1[459]
   PIN dout1[460]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  714.0575 192.83 714.1975 192.97 ;
      END
   END dout1[460]
   PIN dout1[461]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  715.2325 192.83 715.3725 192.97 ;
      END
   END dout1[461]
   PIN dout1[462]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  716.4075 192.83 716.5475 192.97 ;
      END
   END dout1[462]
   PIN dout1[463]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  717.5825 192.83 717.7225 192.97 ;
      END
   END dout1[463]
   PIN dout1[464]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  718.7575 192.83 718.8975 192.97 ;
      END
   END dout1[464]
   PIN dout1[465]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  719.9325 192.83 720.0725 192.97 ;
      END
   END dout1[465]
   PIN dout1[466]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  721.1075 192.83 721.2475 192.97 ;
      END
   END dout1[466]
   PIN dout1[467]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  722.2825 192.83 722.4225 192.97 ;
      END
   END dout1[467]
   PIN dout1[468]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  723.4575 192.83 723.5975 192.97 ;
      END
   END dout1[468]
   PIN dout1[469]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  724.6325 192.83 724.7725 192.97 ;
      END
   END dout1[469]
   PIN dout1[470]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  725.8075 192.83 725.9475 192.97 ;
      END
   END dout1[470]
   PIN dout1[471]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  726.9825 192.83 727.1225 192.97 ;
      END
   END dout1[471]
   PIN dout1[472]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  728.1575 192.83 728.2975 192.97 ;
      END
   END dout1[472]
   PIN dout1[473]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  729.3325 192.83 729.4725 192.97 ;
      END
   END dout1[473]
   PIN dout1[474]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  730.5075 192.83 730.6475 192.97 ;
      END
   END dout1[474]
   PIN dout1[475]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  731.6825 192.83 731.8225 192.97 ;
      END
   END dout1[475]
   PIN dout1[476]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  732.8575 192.83 732.9975 192.97 ;
      END
   END dout1[476]
   PIN dout1[477]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  734.0325 192.83 734.1725 192.97 ;
      END
   END dout1[477]
   PIN dout1[478]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  735.2075 192.83 735.3475 192.97 ;
      END
   END dout1[478]
   PIN dout1[479]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  736.3825 192.83 736.5225 192.97 ;
      END
   END dout1[479]
   PIN dout1[480]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  737.5575 192.83 737.6975 192.97 ;
      END
   END dout1[480]
   PIN dout1[481]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  738.7325 192.83 738.8725 192.97 ;
      END
   END dout1[481]
   PIN dout1[482]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  739.9075 192.83 740.0475 192.97 ;
      END
   END dout1[482]
   PIN dout1[483]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  741.0825 192.83 741.2225 192.97 ;
      END
   END dout1[483]
   PIN dout1[484]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  742.2575 192.83 742.3975 192.97 ;
      END
   END dout1[484]
   PIN dout1[485]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  743.4325 192.83 743.5725 192.97 ;
      END
   END dout1[485]
   PIN dout1[486]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  744.6075 192.83 744.7475 192.97 ;
      END
   END dout1[486]
   PIN dout1[487]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  745.7825 192.83 745.9225 192.97 ;
      END
   END dout1[487]
   PIN dout1[488]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  746.9575 192.83 747.0975 192.97 ;
      END
   END dout1[488]
   PIN dout1[489]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  748.1325 192.83 748.2725 192.97 ;
      END
   END dout1[489]
   PIN dout1[490]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  749.3075 192.83 749.4475 192.97 ;
      END
   END dout1[490]
   PIN dout1[491]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  750.4825 192.83 750.6225 192.97 ;
      END
   END dout1[491]
   PIN dout1[492]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  751.6575 192.83 751.7975 192.97 ;
      END
   END dout1[492]
   PIN dout1[493]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  752.8325 192.83 752.9725 192.97 ;
      END
   END dout1[493]
   PIN dout1[494]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  754.0075 192.83 754.1475 192.97 ;
      END
   END dout1[494]
   PIN dout1[495]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  755.1825 192.83 755.3225 192.97 ;
      END
   END dout1[495]
   PIN dout1[496]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  756.3575 192.83 756.4975 192.97 ;
      END
   END dout1[496]
   PIN dout1[497]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  757.5325 192.83 757.6725 192.97 ;
      END
   END dout1[497]
   PIN dout1[498]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  758.7075 192.83 758.8475 192.97 ;
      END
   END dout1[498]
   PIN dout1[499]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  759.8825 192.83 760.0225 192.97 ;
      END
   END dout1[499]
   PIN dout1[500]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  761.0575 192.83 761.1975 192.97 ;
      END
   END dout1[500]
   PIN dout1[501]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  762.2325 192.83 762.3725 192.97 ;
      END
   END dout1[501]
   PIN dout1[502]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  763.4075 192.83 763.5475 192.97 ;
      END
   END dout1[502]
   PIN dout1[503]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  764.5825 192.83 764.7225 192.97 ;
      END
   END dout1[503]
   PIN dout1[504]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  765.7575 192.83 765.8975 192.97 ;
      END
   END dout1[504]
   PIN dout1[505]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  766.9325 192.83 767.0725 192.97 ;
      END
   END dout1[505]
   PIN dout1[506]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  768.1075 192.83 768.2475 192.97 ;
      END
   END dout1[506]
   PIN dout1[507]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  769.2825 192.83 769.4225 192.97 ;
      END
   END dout1[507]
   PIN dout1[508]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  770.4575 192.83 770.5975 192.97 ;
      END
   END dout1[508]
   PIN dout1[509]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  771.6325 192.83 771.7725 192.97 ;
      END
   END dout1[509]
   PIN dout1[510]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  772.8075 192.83 772.9475 192.97 ;
      END
   END dout1[510]
   PIN dout1[511]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  773.9825 192.83 774.1225 192.97 ;
      END
   END dout1[511]
   PIN dout1[512]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  775.1575 192.83 775.2975 192.97 ;
      END
   END dout1[512]
   PIN dout1[513]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  776.3325 192.83 776.4725 192.97 ;
      END
   END dout1[513]
   PIN dout1[514]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  777.5075 192.83 777.6475 192.97 ;
      END
   END dout1[514]
   PIN dout1[515]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  778.6825 192.83 778.8225 192.97 ;
      END
   END dout1[515]
   PIN dout1[516]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  779.8575 192.83 779.9975 192.97 ;
      END
   END dout1[516]
   PIN dout1[517]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  781.0325 192.83 781.1725 192.97 ;
      END
   END dout1[517]
   PIN dout1[518]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  782.2075 192.83 782.3475 192.97 ;
      END
   END dout1[518]
   PIN dout1[519]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  783.3825 192.83 783.5225 192.97 ;
      END
   END dout1[519]
   PIN dout1[520]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  784.5575 192.83 784.6975 192.97 ;
      END
   END dout1[520]
   PIN dout1[521]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  785.7325 192.83 785.8725 192.97 ;
      END
   END dout1[521]
   PIN dout1[522]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  786.9075 192.83 787.0475 192.97 ;
      END
   END dout1[522]
   PIN dout1[523]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  788.0825 192.83 788.2225 192.97 ;
      END
   END dout1[523]
   PIN dout1[524]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  789.2575 192.83 789.3975 192.97 ;
      END
   END dout1[524]
   PIN dout1[525]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  790.4325 192.83 790.5725 192.97 ;
      END
   END dout1[525]
   PIN dout1[526]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  791.6075 192.83 791.7475 192.97 ;
      END
   END dout1[526]
   PIN dout1[527]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  792.7825 192.83 792.9225 192.97 ;
      END
   END dout1[527]
   PIN dout1[528]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  793.9575 192.83 794.0975 192.97 ;
      END
   END dout1[528]
   PIN dout1[529]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  795.1325 192.83 795.2725 192.97 ;
      END
   END dout1[529]
   PIN dout1[530]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  796.3075 192.83 796.4475 192.97 ;
      END
   END dout1[530]
   PIN dout1[531]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  797.4825 192.83 797.6225 192.97 ;
      END
   END dout1[531]
   PIN dout1[532]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  798.6575 192.83 798.7975 192.97 ;
      END
   END dout1[532]
   PIN dout1[533]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  799.8325 192.83 799.9725 192.97 ;
      END
   END dout1[533]
   PIN dout1[534]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  801.0075 192.83 801.1475 192.97 ;
      END
   END dout1[534]
   PIN dout1[535]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  802.1825 192.83 802.3225 192.97 ;
      END
   END dout1[535]
   PIN dout1[536]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  803.3575 192.83 803.4975 192.97 ;
      END
   END dout1[536]
   PIN dout1[537]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  804.5325 192.83 804.6725 192.97 ;
      END
   END dout1[537]
   PIN dout1[538]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  805.7075 192.83 805.8475 192.97 ;
      END
   END dout1[538]
   PIN dout1[539]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  806.8825 192.83 807.0225 192.97 ;
      END
   END dout1[539]
   PIN dout1[540]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  808.0575 192.83 808.1975 192.97 ;
      END
   END dout1[540]
   PIN dout1[541]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  809.2325 192.83 809.3725 192.97 ;
      END
   END dout1[541]
   PIN dout1[542]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  810.4075 192.83 810.5475 192.97 ;
      END
   END dout1[542]
   PIN dout1[543]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  811.5825 192.83 811.7225 192.97 ;
      END
   END dout1[543]
   PIN dout1[544]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  812.7575 192.83 812.8975 192.97 ;
      END
   END dout1[544]
   PIN dout1[545]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  813.9325 192.83 814.0725 192.97 ;
      END
   END dout1[545]
   PIN dout1[546]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  815.1075 192.83 815.2475 192.97 ;
      END
   END dout1[546]
   PIN dout1[547]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  816.2825 192.83 816.4225 192.97 ;
      END
   END dout1[547]
   PIN dout1[548]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  817.4575 192.83 817.5975 192.97 ;
      END
   END dout1[548]
   PIN dout1[549]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  818.6325 192.83 818.7725 192.97 ;
      END
   END dout1[549]
   PIN dout1[550]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  819.8075 192.83 819.9475 192.97 ;
      END
   END dout1[550]
   PIN dout1[551]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  820.9825 192.83 821.1225 192.97 ;
      END
   END dout1[551]
   PIN dout1[552]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  822.1575 192.83 822.2975 192.97 ;
      END
   END dout1[552]
   PIN dout1[553]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  823.3325 192.83 823.4725 192.97 ;
      END
   END dout1[553]
   PIN dout1[554]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  824.5075 192.83 824.6475 192.97 ;
      END
   END dout1[554]
   PIN dout1[555]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  825.6825 192.83 825.8225 192.97 ;
      END
   END dout1[555]
   PIN dout1[556]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  826.8575 192.83 826.9975 192.97 ;
      END
   END dout1[556]
   PIN dout1[557]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  828.0325 192.83 828.1725 192.97 ;
      END
   END dout1[557]
   PIN dout1[558]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  829.2075 192.83 829.3475 192.97 ;
      END
   END dout1[558]
   PIN dout1[559]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  830.3825 192.83 830.5225 192.97 ;
      END
   END dout1[559]
   PIN dout1[560]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  831.5575 192.83 831.6975 192.97 ;
      END
   END dout1[560]
   PIN dout1[561]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  832.7325 192.83 832.8725 192.97 ;
      END
   END dout1[561]
   PIN dout1[562]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  833.9075 192.83 834.0475 192.97 ;
      END
   END dout1[562]
   PIN dout1[563]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  835.0825 192.83 835.2225 192.97 ;
      END
   END dout1[563]
   PIN dout1[564]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  836.2575 192.83 836.3975 192.97 ;
      END
   END dout1[564]
   PIN dout1[565]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  837.4325 192.83 837.5725 192.97 ;
      END
   END dout1[565]
   PIN dout1[566]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  838.6075 192.83 838.7475 192.97 ;
      END
   END dout1[566]
   PIN dout1[567]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  839.7825 192.83 839.9225 192.97 ;
      END
   END dout1[567]
   PIN dout1[568]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  840.9575 192.83 841.0975 192.97 ;
      END
   END dout1[568]
   PIN dout1[569]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  842.1325 192.83 842.2725 192.97 ;
      END
   END dout1[569]
   PIN dout1[570]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  843.3075 192.83 843.4475 192.97 ;
      END
   END dout1[570]
   PIN dout1[571]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  844.4825 192.83 844.6225 192.97 ;
      END
   END dout1[571]
   PIN dout1[572]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  845.6575 192.83 845.7975 192.97 ;
      END
   END dout1[572]
   PIN dout1[573]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  846.8325 192.83 846.9725 192.97 ;
      END
   END dout1[573]
   PIN dout1[574]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  848.0075 192.83 848.1475 192.97 ;
      END
   END dout1[574]
   PIN dout1[575]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  849.1825 192.83 849.3225 192.97 ;
      END
   END dout1[575]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 1785.15 192.83 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 1785.15 192.83 ;
   LAYER  metal3 ;
      RECT  0.14 0.14 0.28 88.04 ;
      RECT  0.28 0.14 1785.15 88.04 ;
      RECT  0.28 88.04 1785.15 88.46 ;
      RECT  0.28 88.46 1785.15 192.83 ;
      RECT  0.14 88.695 0.28 192.83 ;
   LAYER  metal4 ;
      RECT  0.14 0.14 137.8625 0.42 ;
      RECT  137.8625 0.42 138.5625 192.83 ;
      RECT  138.5625 0.14 140.7225 0.42 ;
      RECT  141.4225 0.14 143.5825 0.42 ;
      RECT  144.2825 0.14 146.4425 0.42 ;
      RECT  147.1425 0.14 149.3025 0.42 ;
      RECT  150.0025 0.14 152.1625 0.42 ;
      RECT  152.8625 0.14 155.0225 0.42 ;
      RECT  155.7225 0.14 157.8825 0.42 ;
      RECT  158.5825 0.14 160.7425 0.42 ;
      RECT  161.4425 0.14 163.6025 0.42 ;
      RECT  164.3025 0.14 166.4625 0.42 ;
      RECT  167.1625 0.14 169.3225 0.42 ;
      RECT  170.0225 0.14 172.1825 0.42 ;
      RECT  172.8825 0.14 175.0425 0.42 ;
      RECT  175.7425 0.14 177.9025 0.42 ;
      RECT  178.6025 0.14 180.7625 0.42 ;
      RECT  181.4625 0.14 183.6225 0.42 ;
      RECT  184.3225 0.14 186.4825 0.42 ;
      RECT  187.1825 0.14 189.3425 0.42 ;
      RECT  190.0425 0.14 192.2025 0.42 ;
      RECT  192.9025 0.14 195.0625 0.42 ;
      RECT  195.7625 0.14 197.9225 0.42 ;
      RECT  198.6225 0.14 200.7825 0.42 ;
      RECT  201.4825 0.14 203.6425 0.42 ;
      RECT  204.3425 0.14 206.5025 0.42 ;
      RECT  207.2025 0.14 209.3625 0.42 ;
      RECT  210.0625 0.14 212.2225 0.42 ;
      RECT  212.9225 0.14 215.0825 0.42 ;
      RECT  215.7825 0.14 217.9425 0.42 ;
      RECT  218.6425 0.14 220.8025 0.42 ;
      RECT  221.5025 0.14 223.6625 0.42 ;
      RECT  224.3625 0.14 226.5225 0.42 ;
      RECT  227.2225 0.14 229.3825 0.42 ;
      RECT  230.0825 0.14 232.2425 0.42 ;
      RECT  232.9425 0.14 235.1025 0.42 ;
      RECT  235.8025 0.14 237.9625 0.42 ;
      RECT  238.6625 0.14 240.8225 0.42 ;
      RECT  241.5225 0.14 243.6825 0.42 ;
      RECT  244.3825 0.14 246.5425 0.42 ;
      RECT  247.2425 0.14 249.4025 0.42 ;
      RECT  250.1025 0.14 252.2625 0.42 ;
      RECT  252.9625 0.14 255.1225 0.42 ;
      RECT  255.8225 0.14 257.9825 0.42 ;
      RECT  258.6825 0.14 260.8425 0.42 ;
      RECT  261.5425 0.14 263.7025 0.42 ;
      RECT  264.4025 0.14 266.5625 0.42 ;
      RECT  267.2625 0.14 269.4225 0.42 ;
      RECT  270.1225 0.14 272.2825 0.42 ;
      RECT  272.9825 0.14 275.1425 0.42 ;
      RECT  275.8425 0.14 278.0025 0.42 ;
      RECT  278.7025 0.14 280.8625 0.42 ;
      RECT  281.5625 0.14 283.7225 0.42 ;
      RECT  284.4225 0.14 286.5825 0.42 ;
      RECT  287.2825 0.14 289.4425 0.42 ;
      RECT  290.1425 0.14 292.3025 0.42 ;
      RECT  293.0025 0.14 295.1625 0.42 ;
      RECT  295.8625 0.14 298.0225 0.42 ;
      RECT  298.7225 0.14 300.8825 0.42 ;
      RECT  301.5825 0.14 303.7425 0.42 ;
      RECT  304.4425 0.14 306.6025 0.42 ;
      RECT  307.3025 0.14 309.4625 0.42 ;
      RECT  310.1625 0.14 312.3225 0.42 ;
      RECT  313.0225 0.14 315.1825 0.42 ;
      RECT  315.8825 0.14 318.0425 0.42 ;
      RECT  318.7425 0.14 320.9025 0.42 ;
      RECT  321.6025 0.14 323.7625 0.42 ;
      RECT  324.4625 0.14 326.6225 0.42 ;
      RECT  327.3225 0.14 329.4825 0.42 ;
      RECT  330.1825 0.14 332.3425 0.42 ;
      RECT  333.0425 0.14 335.2025 0.42 ;
      RECT  335.9025 0.14 338.0625 0.42 ;
      RECT  338.7625 0.14 340.9225 0.42 ;
      RECT  341.6225 0.14 343.7825 0.42 ;
      RECT  344.4825 0.14 346.6425 0.42 ;
      RECT  347.3425 0.14 349.5025 0.42 ;
      RECT  350.2025 0.14 352.3625 0.42 ;
      RECT  353.0625 0.14 355.2225 0.42 ;
      RECT  355.9225 0.14 358.0825 0.42 ;
      RECT  358.7825 0.14 360.9425 0.42 ;
      RECT  361.6425 0.14 363.8025 0.42 ;
      RECT  364.5025 0.14 366.6625 0.42 ;
      RECT  367.3625 0.14 369.5225 0.42 ;
      RECT  370.2225 0.14 372.3825 0.42 ;
      RECT  373.0825 0.14 375.2425 0.42 ;
      RECT  375.9425 0.14 378.1025 0.42 ;
      RECT  378.8025 0.14 380.9625 0.42 ;
      RECT  381.6625 0.14 383.8225 0.42 ;
      RECT  384.5225 0.14 386.6825 0.42 ;
      RECT  387.3825 0.14 389.5425 0.42 ;
      RECT  390.2425 0.14 392.4025 0.42 ;
      RECT  393.1025 0.14 395.2625 0.42 ;
      RECT  395.9625 0.14 398.1225 0.42 ;
      RECT  398.8225 0.14 400.9825 0.42 ;
      RECT  401.6825 0.14 403.8425 0.42 ;
      RECT  404.5425 0.14 406.7025 0.42 ;
      RECT  407.4025 0.14 409.5625 0.42 ;
      RECT  410.2625 0.14 412.4225 0.42 ;
      RECT  413.1225 0.14 415.2825 0.42 ;
      RECT  415.9825 0.14 418.1425 0.42 ;
      RECT  418.8425 0.14 421.0025 0.42 ;
      RECT  421.7025 0.14 423.8625 0.42 ;
      RECT  424.5625 0.14 426.7225 0.42 ;
      RECT  427.4225 0.14 429.5825 0.42 ;
      RECT  430.2825 0.14 432.4425 0.42 ;
      RECT  433.1425 0.14 435.3025 0.42 ;
      RECT  436.0025 0.14 438.1625 0.42 ;
      RECT  438.8625 0.14 441.0225 0.42 ;
      RECT  441.7225 0.14 443.8825 0.42 ;
      RECT  444.5825 0.14 446.7425 0.42 ;
      RECT  447.4425 0.14 449.6025 0.42 ;
      RECT  450.3025 0.14 452.4625 0.42 ;
      RECT  453.1625 0.14 455.3225 0.42 ;
      RECT  456.0225 0.14 458.1825 0.42 ;
      RECT  458.8825 0.14 461.0425 0.42 ;
      RECT  461.7425 0.14 463.9025 0.42 ;
      RECT  464.6025 0.14 466.7625 0.42 ;
      RECT  467.4625 0.14 469.6225 0.42 ;
      RECT  470.3225 0.14 472.4825 0.42 ;
      RECT  473.1825 0.14 475.3425 0.42 ;
      RECT  476.0425 0.14 478.2025 0.42 ;
      RECT  478.9025 0.14 481.0625 0.42 ;
      RECT  481.7625 0.14 483.9225 0.42 ;
      RECT  484.6225 0.14 486.7825 0.42 ;
      RECT  487.4825 0.14 489.6425 0.42 ;
      RECT  490.3425 0.14 492.5025 0.42 ;
      RECT  493.2025 0.14 495.3625 0.42 ;
      RECT  496.0625 0.14 498.2225 0.42 ;
      RECT  498.9225 0.14 501.0825 0.42 ;
      RECT  501.7825 0.14 503.9425 0.42 ;
      RECT  504.6425 0.14 506.8025 0.42 ;
      RECT  507.5025 0.14 509.6625 0.42 ;
      RECT  510.3625 0.14 512.5225 0.42 ;
      RECT  513.2225 0.14 515.3825 0.42 ;
      RECT  516.0825 0.14 518.2425 0.42 ;
      RECT  518.9425 0.14 521.1025 0.42 ;
      RECT  521.8025 0.14 523.9625 0.42 ;
      RECT  524.6625 0.14 526.8225 0.42 ;
      RECT  527.5225 0.14 529.6825 0.42 ;
      RECT  530.3825 0.14 532.5425 0.42 ;
      RECT  533.2425 0.14 535.4025 0.42 ;
      RECT  536.1025 0.14 538.2625 0.42 ;
      RECT  538.9625 0.14 541.1225 0.42 ;
      RECT  541.8225 0.14 543.9825 0.42 ;
      RECT  544.6825 0.14 546.8425 0.42 ;
      RECT  547.5425 0.14 549.7025 0.42 ;
      RECT  550.4025 0.14 552.5625 0.42 ;
      RECT  553.2625 0.14 555.4225 0.42 ;
      RECT  556.1225 0.14 558.2825 0.42 ;
      RECT  558.9825 0.14 561.1425 0.42 ;
      RECT  561.8425 0.14 564.0025 0.42 ;
      RECT  564.7025 0.14 566.8625 0.42 ;
      RECT  567.5625 0.14 569.7225 0.42 ;
      RECT  570.4225 0.14 572.5825 0.42 ;
      RECT  573.2825 0.14 575.4425 0.42 ;
      RECT  576.1425 0.14 578.3025 0.42 ;
      RECT  579.0025 0.14 581.1625 0.42 ;
      RECT  581.8625 0.14 584.0225 0.42 ;
      RECT  584.7225 0.14 586.8825 0.42 ;
      RECT  587.5825 0.14 589.7425 0.42 ;
      RECT  590.4425 0.14 592.6025 0.42 ;
      RECT  593.3025 0.14 595.4625 0.42 ;
      RECT  596.1625 0.14 598.3225 0.42 ;
      RECT  599.0225 0.14 601.1825 0.42 ;
      RECT  601.8825 0.14 604.0425 0.42 ;
      RECT  604.7425 0.14 606.9025 0.42 ;
      RECT  607.6025 0.14 609.7625 0.42 ;
      RECT  610.4625 0.14 612.6225 0.42 ;
      RECT  613.3225 0.14 615.4825 0.42 ;
      RECT  616.1825 0.14 618.3425 0.42 ;
      RECT  619.0425 0.14 621.2025 0.42 ;
      RECT  621.9025 0.14 624.0625 0.42 ;
      RECT  624.7625 0.14 626.9225 0.42 ;
      RECT  627.6225 0.14 629.7825 0.42 ;
      RECT  630.4825 0.14 632.6425 0.42 ;
      RECT  633.3425 0.14 635.5025 0.42 ;
      RECT  636.2025 0.14 638.3625 0.42 ;
      RECT  639.0625 0.14 641.2225 0.42 ;
      RECT  641.9225 0.14 644.0825 0.42 ;
      RECT  644.7825 0.14 646.9425 0.42 ;
      RECT  647.6425 0.14 649.8025 0.42 ;
      RECT  650.5025 0.14 652.6625 0.42 ;
      RECT  653.3625 0.14 655.5225 0.42 ;
      RECT  656.2225 0.14 658.3825 0.42 ;
      RECT  659.0825 0.14 661.2425 0.42 ;
      RECT  661.9425 0.14 664.1025 0.42 ;
      RECT  664.8025 0.14 666.9625 0.42 ;
      RECT  667.6625 0.14 669.8225 0.42 ;
      RECT  670.5225 0.14 672.6825 0.42 ;
      RECT  673.3825 0.14 675.5425 0.42 ;
      RECT  676.2425 0.14 678.4025 0.42 ;
      RECT  679.1025 0.14 681.2625 0.42 ;
      RECT  681.9625 0.14 684.1225 0.42 ;
      RECT  684.8225 0.14 686.9825 0.42 ;
      RECT  687.6825 0.14 689.8425 0.42 ;
      RECT  690.5425 0.14 692.7025 0.42 ;
      RECT  693.4025 0.14 695.5625 0.42 ;
      RECT  696.2625 0.14 698.4225 0.42 ;
      RECT  699.1225 0.14 701.2825 0.42 ;
      RECT  701.9825 0.14 704.1425 0.42 ;
      RECT  704.8425 0.14 707.0025 0.42 ;
      RECT  707.7025 0.14 709.8625 0.42 ;
      RECT  710.5625 0.14 712.7225 0.42 ;
      RECT  713.4225 0.14 715.5825 0.42 ;
      RECT  716.2825 0.14 718.4425 0.42 ;
      RECT  719.1425 0.14 721.3025 0.42 ;
      RECT  722.0025 0.14 724.1625 0.42 ;
      RECT  724.8625 0.14 727.0225 0.42 ;
      RECT  727.7225 0.14 729.8825 0.42 ;
      RECT  730.5825 0.14 732.7425 0.42 ;
      RECT  733.4425 0.14 735.6025 0.42 ;
      RECT  736.3025 0.14 738.4625 0.42 ;
      RECT  739.1625 0.14 741.3225 0.42 ;
      RECT  742.0225 0.14 744.1825 0.42 ;
      RECT  744.8825 0.14 747.0425 0.42 ;
      RECT  747.7425 0.14 749.9025 0.42 ;
      RECT  750.6025 0.14 752.7625 0.42 ;
      RECT  753.4625 0.14 755.6225 0.42 ;
      RECT  756.3225 0.14 758.4825 0.42 ;
      RECT  759.1825 0.14 761.3425 0.42 ;
      RECT  762.0425 0.14 764.2025 0.42 ;
      RECT  764.9025 0.14 767.0625 0.42 ;
      RECT  767.7625 0.14 769.9225 0.42 ;
      RECT  770.6225 0.14 772.7825 0.42 ;
      RECT  773.4825 0.14 775.6425 0.42 ;
      RECT  776.3425 0.14 778.5025 0.42 ;
      RECT  779.2025 0.14 781.3625 0.42 ;
      RECT  782.0625 0.14 784.2225 0.42 ;
      RECT  784.9225 0.14 787.0825 0.42 ;
      RECT  787.7825 0.14 789.9425 0.42 ;
      RECT  790.6425 0.14 792.8025 0.42 ;
      RECT  793.5025 0.14 795.6625 0.42 ;
      RECT  796.3625 0.14 798.5225 0.42 ;
      RECT  799.2225 0.14 801.3825 0.42 ;
      RECT  802.0825 0.14 804.2425 0.42 ;
      RECT  804.9425 0.14 807.1025 0.42 ;
      RECT  807.8025 0.14 809.9625 0.42 ;
      RECT  810.6625 0.14 812.8225 0.42 ;
      RECT  813.5225 0.14 815.6825 0.42 ;
      RECT  816.3825 0.14 818.5425 0.42 ;
      RECT  819.2425 0.14 821.4025 0.42 ;
      RECT  822.1025 0.14 824.2625 0.42 ;
      RECT  824.9625 0.14 827.1225 0.42 ;
      RECT  827.8225 0.14 829.9825 0.42 ;
      RECT  830.6825 0.14 832.8425 0.42 ;
      RECT  833.5425 0.14 835.7025 0.42 ;
      RECT  836.4025 0.14 838.5625 0.42 ;
      RECT  839.2625 0.14 841.4225 0.42 ;
      RECT  842.1225 0.14 844.2825 0.42 ;
      RECT  844.9825 0.14 847.1425 0.42 ;
      RECT  847.8425 0.14 850.0025 0.42 ;
      RECT  850.7025 0.14 852.8625 0.42 ;
      RECT  853.5625 0.14 855.7225 0.42 ;
      RECT  856.4225 0.14 858.5825 0.42 ;
      RECT  859.2825 0.14 861.4425 0.42 ;
      RECT  862.1425 0.14 864.3025 0.42 ;
      RECT  865.0025 0.14 867.1625 0.42 ;
      RECT  867.8625 0.14 870.0225 0.42 ;
      RECT  870.7225 0.14 872.8825 0.42 ;
      RECT  873.5825 0.14 875.7425 0.42 ;
      RECT  876.4425 0.14 878.6025 0.42 ;
      RECT  879.3025 0.14 881.4625 0.42 ;
      RECT  882.1625 0.14 884.3225 0.42 ;
      RECT  885.0225 0.14 887.1825 0.42 ;
      RECT  887.8825 0.14 890.0425 0.42 ;
      RECT  890.7425 0.14 892.9025 0.42 ;
      RECT  893.6025 0.14 895.7625 0.42 ;
      RECT  896.4625 0.14 898.6225 0.42 ;
      RECT  899.3225 0.14 901.4825 0.42 ;
      RECT  902.1825 0.14 904.3425 0.42 ;
      RECT  905.0425 0.14 907.2025 0.42 ;
      RECT  907.9025 0.14 910.0625 0.42 ;
      RECT  910.7625 0.14 912.9225 0.42 ;
      RECT  913.6225 0.14 915.7825 0.42 ;
      RECT  916.4825 0.14 918.6425 0.42 ;
      RECT  919.3425 0.14 921.5025 0.42 ;
      RECT  922.2025 0.14 924.3625 0.42 ;
      RECT  925.0625 0.14 927.2225 0.42 ;
      RECT  927.9225 0.14 930.0825 0.42 ;
      RECT  930.7825 0.14 932.9425 0.42 ;
      RECT  933.6425 0.14 935.8025 0.42 ;
      RECT  936.5025 0.14 938.6625 0.42 ;
      RECT  939.3625 0.14 941.5225 0.42 ;
      RECT  942.2225 0.14 944.3825 0.42 ;
      RECT  945.0825 0.14 947.2425 0.42 ;
      RECT  947.9425 0.14 950.1025 0.42 ;
      RECT  950.8025 0.14 952.9625 0.42 ;
      RECT  953.6625 0.14 955.8225 0.42 ;
      RECT  956.5225 0.14 958.6825 0.42 ;
      RECT  959.3825 0.14 961.5425 0.42 ;
      RECT  962.2425 0.14 964.4025 0.42 ;
      RECT  965.1025 0.14 967.2625 0.42 ;
      RECT  967.9625 0.14 970.1225 0.42 ;
      RECT  970.8225 0.14 972.9825 0.42 ;
      RECT  973.6825 0.14 975.8425 0.42 ;
      RECT  976.5425 0.14 978.7025 0.42 ;
      RECT  979.4025 0.14 981.5625 0.42 ;
      RECT  982.2625 0.14 984.4225 0.42 ;
      RECT  985.1225 0.14 987.2825 0.42 ;
      RECT  987.9825 0.14 990.1425 0.42 ;
      RECT  990.8425 0.14 993.0025 0.42 ;
      RECT  993.7025 0.14 995.8625 0.42 ;
      RECT  996.5625 0.14 998.7225 0.42 ;
      RECT  999.4225 0.14 1001.5825 0.42 ;
      RECT  1002.2825 0.14 1004.4425 0.42 ;
      RECT  1005.1425 0.14 1007.3025 0.42 ;
      RECT  1008.0025 0.14 1010.1625 0.42 ;
      RECT  1010.8625 0.14 1013.0225 0.42 ;
      RECT  1013.7225 0.14 1015.8825 0.42 ;
      RECT  1016.5825 0.14 1018.7425 0.42 ;
      RECT  1019.4425 0.14 1021.6025 0.42 ;
      RECT  1022.3025 0.14 1024.4625 0.42 ;
      RECT  1025.1625 0.14 1027.3225 0.42 ;
      RECT  1028.0225 0.14 1030.1825 0.42 ;
      RECT  1030.8825 0.14 1033.0425 0.42 ;
      RECT  1033.7425 0.14 1035.9025 0.42 ;
      RECT  1036.6025 0.14 1038.7625 0.42 ;
      RECT  1039.4625 0.14 1041.6225 0.42 ;
      RECT  1042.3225 0.14 1044.4825 0.42 ;
      RECT  1045.1825 0.14 1047.3425 0.42 ;
      RECT  1048.0425 0.14 1050.2025 0.42 ;
      RECT  1050.9025 0.14 1053.0625 0.42 ;
      RECT  1053.7625 0.14 1055.9225 0.42 ;
      RECT  1056.6225 0.14 1058.7825 0.42 ;
      RECT  1059.4825 0.14 1061.6425 0.42 ;
      RECT  1062.3425 0.14 1064.5025 0.42 ;
      RECT  1065.2025 0.14 1067.3625 0.42 ;
      RECT  1068.0625 0.14 1070.2225 0.42 ;
      RECT  1070.9225 0.14 1073.0825 0.42 ;
      RECT  1073.7825 0.14 1075.9425 0.42 ;
      RECT  1076.6425 0.14 1078.8025 0.42 ;
      RECT  1079.5025 0.14 1081.6625 0.42 ;
      RECT  1082.3625 0.14 1084.5225 0.42 ;
      RECT  1085.2225 0.14 1087.3825 0.42 ;
      RECT  1088.0825 0.14 1090.2425 0.42 ;
      RECT  1090.9425 0.14 1093.1025 0.42 ;
      RECT  1093.8025 0.14 1095.9625 0.42 ;
      RECT  1096.6625 0.14 1098.8225 0.42 ;
      RECT  1099.5225 0.14 1101.6825 0.42 ;
      RECT  1102.3825 0.14 1104.5425 0.42 ;
      RECT  1105.2425 0.14 1107.4025 0.42 ;
      RECT  1108.1025 0.14 1110.2625 0.42 ;
      RECT  1110.9625 0.14 1113.1225 0.42 ;
      RECT  1113.8225 0.14 1115.9825 0.42 ;
      RECT  1116.6825 0.14 1118.8425 0.42 ;
      RECT  1119.5425 0.14 1121.7025 0.42 ;
      RECT  1122.4025 0.14 1124.5625 0.42 ;
      RECT  1125.2625 0.14 1127.4225 0.42 ;
      RECT  1128.1225 0.14 1130.2825 0.42 ;
      RECT  1130.9825 0.14 1133.1425 0.42 ;
      RECT  1133.8425 0.14 1136.0025 0.42 ;
      RECT  1136.7025 0.14 1138.8625 0.42 ;
      RECT  1139.5625 0.14 1141.7225 0.42 ;
      RECT  1142.4225 0.14 1144.5825 0.42 ;
      RECT  1145.2825 0.14 1147.4425 0.42 ;
      RECT  1148.1425 0.14 1150.3025 0.42 ;
      RECT  1151.0025 0.14 1153.1625 0.42 ;
      RECT  1153.8625 0.14 1156.0225 0.42 ;
      RECT  1156.7225 0.14 1158.8825 0.42 ;
      RECT  1159.5825 0.14 1161.7425 0.42 ;
      RECT  1162.4425 0.14 1164.6025 0.42 ;
      RECT  1165.3025 0.14 1167.4625 0.42 ;
      RECT  1168.1625 0.14 1170.3225 0.42 ;
      RECT  1171.0225 0.14 1173.1825 0.42 ;
      RECT  1173.8825 0.14 1176.0425 0.42 ;
      RECT  1176.7425 0.14 1178.9025 0.42 ;
      RECT  1179.6025 0.14 1181.7625 0.42 ;
      RECT  1182.4625 0.14 1184.6225 0.42 ;
      RECT  1185.3225 0.14 1187.4825 0.42 ;
      RECT  1188.1825 0.14 1190.3425 0.42 ;
      RECT  1191.0425 0.14 1193.2025 0.42 ;
      RECT  1193.9025 0.14 1196.0625 0.42 ;
      RECT  1196.7625 0.14 1198.9225 0.42 ;
      RECT  1199.6225 0.14 1201.7825 0.42 ;
      RECT  1202.4825 0.14 1204.6425 0.42 ;
      RECT  1205.3425 0.14 1207.5025 0.42 ;
      RECT  1208.2025 0.14 1210.3625 0.42 ;
      RECT  1211.0625 0.14 1213.2225 0.42 ;
      RECT  1213.9225 0.14 1216.0825 0.42 ;
      RECT  1216.7825 0.14 1218.9425 0.42 ;
      RECT  1219.6425 0.14 1221.8025 0.42 ;
      RECT  1222.5025 0.14 1224.6625 0.42 ;
      RECT  1225.3625 0.14 1227.5225 0.42 ;
      RECT  1228.2225 0.14 1230.3825 0.42 ;
      RECT  1231.0825 0.14 1233.2425 0.42 ;
      RECT  1233.9425 0.14 1236.1025 0.42 ;
      RECT  1236.8025 0.14 1238.9625 0.42 ;
      RECT  1239.6625 0.14 1241.8225 0.42 ;
      RECT  1242.5225 0.14 1244.6825 0.42 ;
      RECT  1245.3825 0.14 1247.5425 0.42 ;
      RECT  1248.2425 0.14 1250.4025 0.42 ;
      RECT  1251.1025 0.14 1253.2625 0.42 ;
      RECT  1253.9625 0.14 1256.1225 0.42 ;
      RECT  1256.8225 0.14 1258.9825 0.42 ;
      RECT  1259.6825 0.14 1261.8425 0.42 ;
      RECT  1262.5425 0.14 1264.7025 0.42 ;
      RECT  1265.4025 0.14 1267.5625 0.42 ;
      RECT  1268.2625 0.14 1270.4225 0.42 ;
      RECT  1271.1225 0.14 1273.2825 0.42 ;
      RECT  1273.9825 0.14 1276.1425 0.42 ;
      RECT  1276.8425 0.14 1279.0025 0.42 ;
      RECT  1279.7025 0.14 1281.8625 0.42 ;
      RECT  1282.5625 0.14 1284.7225 0.42 ;
      RECT  1285.4225 0.14 1287.5825 0.42 ;
      RECT  1288.2825 0.14 1290.4425 0.42 ;
      RECT  1291.1425 0.14 1293.3025 0.42 ;
      RECT  1294.0025 0.14 1296.1625 0.42 ;
      RECT  1296.8625 0.14 1299.0225 0.42 ;
      RECT  1299.7225 0.14 1301.8825 0.42 ;
      RECT  1302.5825 0.14 1304.7425 0.42 ;
      RECT  1305.4425 0.14 1307.6025 0.42 ;
      RECT  1308.3025 0.14 1310.4625 0.42 ;
      RECT  1311.1625 0.14 1313.3225 0.42 ;
      RECT  1314.0225 0.14 1316.1825 0.42 ;
      RECT  1316.8825 0.14 1319.0425 0.42 ;
      RECT  1319.7425 0.14 1321.9025 0.42 ;
      RECT  1322.6025 0.14 1324.7625 0.42 ;
      RECT  1325.4625 0.14 1327.6225 0.42 ;
      RECT  1328.3225 0.14 1330.4825 0.42 ;
      RECT  1331.1825 0.14 1333.3425 0.42 ;
      RECT  1334.0425 0.14 1336.2025 0.42 ;
      RECT  1336.9025 0.14 1339.0625 0.42 ;
      RECT  1339.7625 0.14 1341.9225 0.42 ;
      RECT  1342.6225 0.14 1344.7825 0.42 ;
      RECT  1345.4825 0.14 1347.6425 0.42 ;
      RECT  1348.3425 0.14 1350.5025 0.42 ;
      RECT  1351.2025 0.14 1353.3625 0.42 ;
      RECT  1354.0625 0.14 1356.2225 0.42 ;
      RECT  1356.9225 0.14 1359.0825 0.42 ;
      RECT  1359.7825 0.14 1361.9425 0.42 ;
      RECT  1362.6425 0.14 1364.8025 0.42 ;
      RECT  1365.5025 0.14 1367.6625 0.42 ;
      RECT  1368.3625 0.14 1370.5225 0.42 ;
      RECT  1371.2225 0.14 1373.3825 0.42 ;
      RECT  1374.0825 0.14 1376.2425 0.42 ;
      RECT  1376.9425 0.14 1379.1025 0.42 ;
      RECT  1379.8025 0.14 1381.9625 0.42 ;
      RECT  1382.6625 0.14 1384.8225 0.42 ;
      RECT  1385.5225 0.14 1387.6825 0.42 ;
      RECT  1388.3825 0.14 1390.5425 0.42 ;
      RECT  1391.2425 0.14 1393.4025 0.42 ;
      RECT  1394.1025 0.14 1396.2625 0.42 ;
      RECT  1396.9625 0.14 1399.1225 0.42 ;
      RECT  1399.8225 0.14 1401.9825 0.42 ;
      RECT  1402.6825 0.14 1404.8425 0.42 ;
      RECT  1405.5425 0.14 1407.7025 0.42 ;
      RECT  1408.4025 0.14 1410.5625 0.42 ;
      RECT  1411.2625 0.14 1413.4225 0.42 ;
      RECT  1414.1225 0.14 1416.2825 0.42 ;
      RECT  1416.9825 0.14 1419.1425 0.42 ;
      RECT  1419.8425 0.14 1422.0025 0.42 ;
      RECT  1422.7025 0.14 1424.8625 0.42 ;
      RECT  1425.5625 0.14 1427.7225 0.42 ;
      RECT  1428.4225 0.14 1430.5825 0.42 ;
      RECT  1431.2825 0.14 1433.4425 0.42 ;
      RECT  1434.1425 0.14 1436.3025 0.42 ;
      RECT  1437.0025 0.14 1439.1625 0.42 ;
      RECT  1439.8625 0.14 1442.0225 0.42 ;
      RECT  1442.7225 0.14 1444.8825 0.42 ;
      RECT  1445.5825 0.14 1447.7425 0.42 ;
      RECT  1448.4425 0.14 1450.6025 0.42 ;
      RECT  1451.3025 0.14 1453.4625 0.42 ;
      RECT  1454.1625 0.14 1456.3225 0.42 ;
      RECT  1457.0225 0.14 1459.1825 0.42 ;
      RECT  1459.8825 0.14 1462.0425 0.42 ;
      RECT  1462.7425 0.14 1464.9025 0.42 ;
      RECT  1465.6025 0.14 1467.7625 0.42 ;
      RECT  1468.4625 0.14 1470.6225 0.42 ;
      RECT  1471.3225 0.14 1473.4825 0.42 ;
      RECT  1474.1825 0.14 1476.3425 0.42 ;
      RECT  1477.0425 0.14 1479.2025 0.42 ;
      RECT  1479.9025 0.14 1482.0625 0.42 ;
      RECT  1482.7625 0.14 1484.9225 0.42 ;
      RECT  1485.6225 0.14 1487.7825 0.42 ;
      RECT  1488.4825 0.14 1490.6425 0.42 ;
      RECT  1491.3425 0.14 1493.5025 0.42 ;
      RECT  1494.2025 0.14 1496.3625 0.42 ;
      RECT  1497.0625 0.14 1499.2225 0.42 ;
      RECT  1499.9225 0.14 1502.0825 0.42 ;
      RECT  1502.7825 0.14 1504.9425 0.42 ;
      RECT  1505.6425 0.14 1507.8025 0.42 ;
      RECT  1508.5025 0.14 1510.6625 0.42 ;
      RECT  1511.3625 0.14 1513.5225 0.42 ;
      RECT  1514.2225 0.14 1516.3825 0.42 ;
      RECT  1517.0825 0.14 1519.2425 0.42 ;
      RECT  1519.9425 0.14 1522.1025 0.42 ;
      RECT  1522.8025 0.14 1524.9625 0.42 ;
      RECT  1525.6625 0.14 1527.8225 0.42 ;
      RECT  1528.5225 0.14 1530.6825 0.42 ;
      RECT  1531.3825 0.14 1533.5425 0.42 ;
      RECT  1534.2425 0.14 1536.4025 0.42 ;
      RECT  1537.1025 0.14 1539.2625 0.42 ;
      RECT  1539.9625 0.14 1542.1225 0.42 ;
      RECT  1542.8225 0.14 1544.9825 0.42 ;
      RECT  1545.6825 0.14 1547.8425 0.42 ;
      RECT  1548.5425 0.14 1550.7025 0.42 ;
      RECT  1551.4025 0.14 1553.5625 0.42 ;
      RECT  1554.2625 0.14 1556.4225 0.42 ;
      RECT  1557.1225 0.14 1559.2825 0.42 ;
      RECT  1559.9825 0.14 1562.1425 0.42 ;
      RECT  1562.8425 0.14 1565.0025 0.42 ;
      RECT  1565.7025 0.14 1567.8625 0.42 ;
      RECT  1568.5625 0.14 1570.7225 0.42 ;
      RECT  1571.4225 0.14 1573.5825 0.42 ;
      RECT  1574.2825 0.14 1576.4425 0.42 ;
      RECT  1577.1425 0.14 1579.3025 0.42 ;
      RECT  1580.0025 0.14 1582.1625 0.42 ;
      RECT  1582.8625 0.14 1585.0225 0.42 ;
      RECT  1585.7225 0.14 1587.8825 0.42 ;
      RECT  1588.5825 0.14 1590.7425 0.42 ;
      RECT  1591.4425 0.14 1593.6025 0.42 ;
      RECT  1594.3025 0.14 1596.4625 0.42 ;
      RECT  1597.1625 0.14 1599.3225 0.42 ;
      RECT  1600.0225 0.14 1602.1825 0.42 ;
      RECT  1602.8825 0.14 1605.0425 0.42 ;
      RECT  1605.7425 0.14 1607.9025 0.42 ;
      RECT  1608.6025 0.14 1610.7625 0.42 ;
      RECT  1611.4625 0.14 1613.6225 0.42 ;
      RECT  1614.3225 0.14 1616.4825 0.42 ;
      RECT  1617.1825 0.14 1619.3425 0.42 ;
      RECT  1620.0425 0.14 1622.2025 0.42 ;
      RECT  1622.9025 0.14 1625.0625 0.42 ;
      RECT  1625.7625 0.14 1627.9225 0.42 ;
      RECT  1628.6225 0.14 1630.7825 0.42 ;
      RECT  1631.4825 0.14 1633.6425 0.42 ;
      RECT  1634.3425 0.14 1636.5025 0.42 ;
      RECT  1637.2025 0.14 1639.3625 0.42 ;
      RECT  1640.0625 0.14 1642.2225 0.42 ;
      RECT  1642.9225 0.14 1645.0825 0.42 ;
      RECT  1645.7825 0.14 1647.9425 0.42 ;
      RECT  1648.6425 0.14 1650.8025 0.42 ;
      RECT  1651.5025 0.14 1653.6625 0.42 ;
      RECT  1654.3625 0.14 1656.5225 0.42 ;
      RECT  1657.2225 0.14 1659.3825 0.42 ;
      RECT  1660.0825 0.14 1662.2425 0.42 ;
      RECT  1662.9425 0.14 1665.1025 0.42 ;
      RECT  1665.8025 0.14 1667.9625 0.42 ;
      RECT  1668.6625 0.14 1670.8225 0.42 ;
      RECT  1671.5225 0.14 1673.6825 0.42 ;
      RECT  1674.3825 0.14 1676.5425 0.42 ;
      RECT  1677.2425 0.14 1679.4025 0.42 ;
      RECT  1680.1025 0.14 1682.2625 0.42 ;
      RECT  1682.9625 0.14 1685.1225 0.42 ;
      RECT  1685.8225 0.14 1687.9825 0.42 ;
      RECT  1688.6825 0.14 1690.8425 0.42 ;
      RECT  1691.5425 0.14 1693.7025 0.42 ;
      RECT  1694.4025 0.14 1696.5625 0.42 ;
      RECT  1697.2625 0.14 1699.4225 0.42 ;
      RECT  1700.1225 0.14 1702.2825 0.42 ;
      RECT  1702.9825 0.14 1705.1425 0.42 ;
      RECT  1705.8425 0.14 1708.0025 0.42 ;
      RECT  1708.7025 0.14 1710.8625 0.42 ;
      RECT  1711.5625 0.14 1713.7225 0.42 ;
      RECT  1714.4225 0.14 1716.5825 0.42 ;
      RECT  1717.2825 0.14 1719.4425 0.42 ;
      RECT  1720.1425 0.14 1722.3025 0.42 ;
      RECT  1723.0025 0.14 1725.1625 0.42 ;
      RECT  1725.8625 0.14 1728.0225 0.42 ;
      RECT  1728.7225 0.14 1730.8825 0.42 ;
      RECT  1731.5825 0.14 1733.7425 0.42 ;
      RECT  1734.4425 0.14 1736.6025 0.42 ;
      RECT  1737.3025 0.14 1739.4625 0.42 ;
      RECT  1740.1625 0.14 1742.3225 0.42 ;
      RECT  1743.0225 0.14 1745.1825 0.42 ;
      RECT  1745.8825 0.14 1748.0425 0.42 ;
      RECT  1748.7425 0.14 1750.9025 0.42 ;
      RECT  1751.6025 0.14 1753.7625 0.42 ;
      RECT  1754.4625 0.14 1756.6225 0.42 ;
      RECT  1757.3225 0.14 1759.4825 0.42 ;
      RECT  1760.1825 0.14 1762.3425 0.42 ;
      RECT  1763.0425 0.14 1765.2025 0.42 ;
      RECT  1765.9025 0.14 1768.0625 0.42 ;
      RECT  1768.7625 0.14 1770.9225 0.42 ;
      RECT  1771.6225 0.14 1773.7825 0.42 ;
      RECT  1774.4825 0.14 1776.6425 0.42 ;
      RECT  1777.3425 0.14 1779.5025 0.42 ;
      RECT  1780.2025 0.14 1782.3625 0.42 ;
      RECT  1783.0625 0.14 1785.15 0.42 ;
      RECT  0.14 0.42 132.715 192.55 ;
      RECT  132.715 0.42 133.415 192.55 ;
      RECT  133.415 0.42 137.8625 192.55 ;
      RECT  133.415 192.55 137.8625 192.83 ;
      RECT  0.14 192.55 131.575 192.83 ;
      RECT  138.5625 0.42 891.35 192.55 ;
      RECT  891.35 0.42 892.05 192.55 ;
      RECT  892.05 0.42 1785.15 192.55 ;
      RECT  1021.1125 192.55 1785.15 192.83 ;
      RECT  892.62 192.55 1014.215 192.83 ;
      RECT  1014.915 192.55 1020.4125 192.83 ;
      RECT  138.5625 192.55 173.2775 192.83 ;
      RECT  173.9775 192.55 174.4525 192.83 ;
      RECT  175.1525 192.55 175.6275 192.83 ;
      RECT  176.3275 192.55 176.8025 192.83 ;
      RECT  177.5025 192.55 177.9775 192.83 ;
      RECT  178.6775 192.55 179.1525 192.83 ;
      RECT  179.8525 192.55 180.3275 192.83 ;
      RECT  181.0275 192.55 181.5025 192.83 ;
      RECT  182.2025 192.55 182.6775 192.83 ;
      RECT  183.3775 192.55 183.8525 192.83 ;
      RECT  184.5525 192.55 185.0275 192.83 ;
      RECT  185.7275 192.55 186.2025 192.83 ;
      RECT  186.9025 192.55 187.3775 192.83 ;
      RECT  188.0775 192.55 188.5525 192.83 ;
      RECT  189.2525 192.55 189.7275 192.83 ;
      RECT  190.4275 192.55 190.9025 192.83 ;
      RECT  191.6025 192.55 192.0775 192.83 ;
      RECT  192.7775 192.55 193.2525 192.83 ;
      RECT  193.9525 192.55 194.4275 192.83 ;
      RECT  195.1275 192.55 195.6025 192.83 ;
      RECT  196.3025 192.55 196.7775 192.83 ;
      RECT  197.4775 192.55 197.9525 192.83 ;
      RECT  198.6525 192.55 199.1275 192.83 ;
      RECT  199.8275 192.55 200.3025 192.83 ;
      RECT  201.0025 192.55 201.4775 192.83 ;
      RECT  202.1775 192.55 202.6525 192.83 ;
      RECT  203.3525 192.55 203.8275 192.83 ;
      RECT  204.5275 192.55 205.0025 192.83 ;
      RECT  205.7025 192.55 206.1775 192.83 ;
      RECT  206.8775 192.55 207.3525 192.83 ;
      RECT  208.0525 192.55 208.5275 192.83 ;
      RECT  209.2275 192.55 209.7025 192.83 ;
      RECT  210.4025 192.55 210.8775 192.83 ;
      RECT  211.5775 192.55 212.0525 192.83 ;
      RECT  212.7525 192.55 213.2275 192.83 ;
      RECT  213.9275 192.55 214.4025 192.83 ;
      RECT  215.1025 192.55 215.5775 192.83 ;
      RECT  216.2775 192.55 216.7525 192.83 ;
      RECT  217.4525 192.55 217.9275 192.83 ;
      RECT  218.6275 192.55 219.1025 192.83 ;
      RECT  219.8025 192.55 220.2775 192.83 ;
      RECT  220.9775 192.55 221.4525 192.83 ;
      RECT  222.1525 192.55 222.6275 192.83 ;
      RECT  223.3275 192.55 223.8025 192.83 ;
      RECT  224.5025 192.55 224.9775 192.83 ;
      RECT  225.6775 192.55 226.1525 192.83 ;
      RECT  226.8525 192.55 227.3275 192.83 ;
      RECT  228.0275 192.55 228.5025 192.83 ;
      RECT  229.2025 192.55 229.6775 192.83 ;
      RECT  230.3775 192.55 230.8525 192.83 ;
      RECT  231.5525 192.55 232.0275 192.83 ;
      RECT  232.7275 192.55 233.2025 192.83 ;
      RECT  233.9025 192.55 234.3775 192.83 ;
      RECT  235.0775 192.55 235.5525 192.83 ;
      RECT  236.2525 192.55 236.7275 192.83 ;
      RECT  237.4275 192.55 237.9025 192.83 ;
      RECT  238.6025 192.55 239.0775 192.83 ;
      RECT  239.7775 192.55 240.2525 192.83 ;
      RECT  240.9525 192.55 241.4275 192.83 ;
      RECT  242.1275 192.55 242.6025 192.83 ;
      RECT  243.3025 192.55 243.7775 192.83 ;
      RECT  244.4775 192.55 244.9525 192.83 ;
      RECT  245.6525 192.55 246.1275 192.83 ;
      RECT  246.8275 192.55 247.3025 192.83 ;
      RECT  248.0025 192.55 248.4775 192.83 ;
      RECT  249.1775 192.55 249.6525 192.83 ;
      RECT  250.3525 192.55 250.8275 192.83 ;
      RECT  251.5275 192.55 252.0025 192.83 ;
      RECT  252.7025 192.55 253.1775 192.83 ;
      RECT  253.8775 192.55 254.3525 192.83 ;
      RECT  255.0525 192.55 255.5275 192.83 ;
      RECT  256.2275 192.55 256.7025 192.83 ;
      RECT  257.4025 192.55 257.8775 192.83 ;
      RECT  258.5775 192.55 259.0525 192.83 ;
      RECT  259.7525 192.55 260.2275 192.83 ;
      RECT  260.9275 192.55 261.4025 192.83 ;
      RECT  262.1025 192.55 262.5775 192.83 ;
      RECT  263.2775 192.55 263.7525 192.83 ;
      RECT  264.4525 192.55 264.9275 192.83 ;
      RECT  265.6275 192.55 266.1025 192.83 ;
      RECT  266.8025 192.55 267.2775 192.83 ;
      RECT  267.9775 192.55 268.4525 192.83 ;
      RECT  269.1525 192.55 269.6275 192.83 ;
      RECT  270.3275 192.55 270.8025 192.83 ;
      RECT  271.5025 192.55 271.9775 192.83 ;
      RECT  272.6775 192.55 273.1525 192.83 ;
      RECT  273.8525 192.55 274.3275 192.83 ;
      RECT  275.0275 192.55 275.5025 192.83 ;
      RECT  276.2025 192.55 276.6775 192.83 ;
      RECT  277.3775 192.55 277.8525 192.83 ;
      RECT  278.5525 192.55 279.0275 192.83 ;
      RECT  279.7275 192.55 280.2025 192.83 ;
      RECT  280.9025 192.55 281.3775 192.83 ;
      RECT  282.0775 192.55 282.5525 192.83 ;
      RECT  283.2525 192.55 283.7275 192.83 ;
      RECT  284.4275 192.55 284.9025 192.83 ;
      RECT  285.6025 192.55 286.0775 192.83 ;
      RECT  286.7775 192.55 287.2525 192.83 ;
      RECT  287.9525 192.55 288.4275 192.83 ;
      RECT  289.1275 192.55 289.6025 192.83 ;
      RECT  290.3025 192.55 290.7775 192.83 ;
      RECT  291.4775 192.55 291.9525 192.83 ;
      RECT  292.6525 192.55 293.1275 192.83 ;
      RECT  293.8275 192.55 294.3025 192.83 ;
      RECT  295.0025 192.55 295.4775 192.83 ;
      RECT  296.1775 192.55 296.6525 192.83 ;
      RECT  297.3525 192.55 297.8275 192.83 ;
      RECT  298.5275 192.55 299.0025 192.83 ;
      RECT  299.7025 192.55 300.1775 192.83 ;
      RECT  300.8775 192.55 301.3525 192.83 ;
      RECT  302.0525 192.55 302.5275 192.83 ;
      RECT  303.2275 192.55 303.7025 192.83 ;
      RECT  304.4025 192.55 304.8775 192.83 ;
      RECT  305.5775 192.55 306.0525 192.83 ;
      RECT  306.7525 192.55 307.2275 192.83 ;
      RECT  307.9275 192.55 308.4025 192.83 ;
      RECT  309.1025 192.55 309.5775 192.83 ;
      RECT  310.2775 192.55 310.7525 192.83 ;
      RECT  311.4525 192.55 311.9275 192.83 ;
      RECT  312.6275 192.55 313.1025 192.83 ;
      RECT  313.8025 192.55 314.2775 192.83 ;
      RECT  314.9775 192.55 315.4525 192.83 ;
      RECT  316.1525 192.55 316.6275 192.83 ;
      RECT  317.3275 192.55 317.8025 192.83 ;
      RECT  318.5025 192.55 318.9775 192.83 ;
      RECT  319.6775 192.55 320.1525 192.83 ;
      RECT  320.8525 192.55 321.3275 192.83 ;
      RECT  322.0275 192.55 322.5025 192.83 ;
      RECT  323.2025 192.55 323.6775 192.83 ;
      RECT  324.3775 192.55 324.8525 192.83 ;
      RECT  325.5525 192.55 326.0275 192.83 ;
      RECT  326.7275 192.55 327.2025 192.83 ;
      RECT  327.9025 192.55 328.3775 192.83 ;
      RECT  329.0775 192.55 329.5525 192.83 ;
      RECT  330.2525 192.55 330.7275 192.83 ;
      RECT  331.4275 192.55 331.9025 192.83 ;
      RECT  332.6025 192.55 333.0775 192.83 ;
      RECT  333.7775 192.55 334.2525 192.83 ;
      RECT  334.9525 192.55 335.4275 192.83 ;
      RECT  336.1275 192.55 336.6025 192.83 ;
      RECT  337.3025 192.55 337.7775 192.83 ;
      RECT  338.4775 192.55 338.9525 192.83 ;
      RECT  339.6525 192.55 340.1275 192.83 ;
      RECT  340.8275 192.55 341.3025 192.83 ;
      RECT  342.0025 192.55 342.4775 192.83 ;
      RECT  343.1775 192.55 343.6525 192.83 ;
      RECT  344.3525 192.55 344.8275 192.83 ;
      RECT  345.5275 192.55 346.0025 192.83 ;
      RECT  346.7025 192.55 347.1775 192.83 ;
      RECT  347.8775 192.55 348.3525 192.83 ;
      RECT  349.0525 192.55 349.5275 192.83 ;
      RECT  350.2275 192.55 350.7025 192.83 ;
      RECT  351.4025 192.55 351.8775 192.83 ;
      RECT  352.5775 192.55 353.0525 192.83 ;
      RECT  353.7525 192.55 354.2275 192.83 ;
      RECT  354.9275 192.55 355.4025 192.83 ;
      RECT  356.1025 192.55 356.5775 192.83 ;
      RECT  357.2775 192.55 357.7525 192.83 ;
      RECT  358.4525 192.55 358.9275 192.83 ;
      RECT  359.6275 192.55 360.1025 192.83 ;
      RECT  360.8025 192.55 361.2775 192.83 ;
      RECT  361.9775 192.55 362.4525 192.83 ;
      RECT  363.1525 192.55 363.6275 192.83 ;
      RECT  364.3275 192.55 364.8025 192.83 ;
      RECT  365.5025 192.55 365.9775 192.83 ;
      RECT  366.6775 192.55 367.1525 192.83 ;
      RECT  367.8525 192.55 368.3275 192.83 ;
      RECT  369.0275 192.55 369.5025 192.83 ;
      RECT  370.2025 192.55 370.6775 192.83 ;
      RECT  371.3775 192.55 371.8525 192.83 ;
      RECT  372.5525 192.55 373.0275 192.83 ;
      RECT  373.7275 192.55 374.2025 192.83 ;
      RECT  374.9025 192.55 375.3775 192.83 ;
      RECT  376.0775 192.55 376.5525 192.83 ;
      RECT  377.2525 192.55 377.7275 192.83 ;
      RECT  378.4275 192.55 378.9025 192.83 ;
      RECT  379.6025 192.55 380.0775 192.83 ;
      RECT  380.7775 192.55 381.2525 192.83 ;
      RECT  381.9525 192.55 382.4275 192.83 ;
      RECT  383.1275 192.55 383.6025 192.83 ;
      RECT  384.3025 192.55 384.7775 192.83 ;
      RECT  385.4775 192.55 385.9525 192.83 ;
      RECT  386.6525 192.55 387.1275 192.83 ;
      RECT  387.8275 192.55 388.3025 192.83 ;
      RECT  389.0025 192.55 389.4775 192.83 ;
      RECT  390.1775 192.55 390.6525 192.83 ;
      RECT  391.3525 192.55 391.8275 192.83 ;
      RECT  392.5275 192.55 393.0025 192.83 ;
      RECT  393.7025 192.55 394.1775 192.83 ;
      RECT  394.8775 192.55 395.3525 192.83 ;
      RECT  396.0525 192.55 396.5275 192.83 ;
      RECT  397.2275 192.55 397.7025 192.83 ;
      RECT  398.4025 192.55 398.8775 192.83 ;
      RECT  399.5775 192.55 400.0525 192.83 ;
      RECT  400.7525 192.55 401.2275 192.83 ;
      RECT  401.9275 192.55 402.4025 192.83 ;
      RECT  403.1025 192.55 403.5775 192.83 ;
      RECT  404.2775 192.55 404.7525 192.83 ;
      RECT  405.4525 192.55 405.9275 192.83 ;
      RECT  406.6275 192.55 407.1025 192.83 ;
      RECT  407.8025 192.55 408.2775 192.83 ;
      RECT  408.9775 192.55 409.4525 192.83 ;
      RECT  410.1525 192.55 410.6275 192.83 ;
      RECT  411.3275 192.55 411.8025 192.83 ;
      RECT  412.5025 192.55 412.9775 192.83 ;
      RECT  413.6775 192.55 414.1525 192.83 ;
      RECT  414.8525 192.55 415.3275 192.83 ;
      RECT  416.0275 192.55 416.5025 192.83 ;
      RECT  417.2025 192.55 417.6775 192.83 ;
      RECT  418.3775 192.55 418.8525 192.83 ;
      RECT  419.5525 192.55 420.0275 192.83 ;
      RECT  420.7275 192.55 421.2025 192.83 ;
      RECT  421.9025 192.55 422.3775 192.83 ;
      RECT  423.0775 192.55 423.5525 192.83 ;
      RECT  424.2525 192.55 424.7275 192.83 ;
      RECT  425.4275 192.55 425.9025 192.83 ;
      RECT  426.6025 192.55 427.0775 192.83 ;
      RECT  427.7775 192.55 428.2525 192.83 ;
      RECT  428.9525 192.55 429.4275 192.83 ;
      RECT  430.1275 192.55 430.6025 192.83 ;
      RECT  431.3025 192.55 431.7775 192.83 ;
      RECT  432.4775 192.55 432.9525 192.83 ;
      RECT  433.6525 192.55 434.1275 192.83 ;
      RECT  434.8275 192.55 435.3025 192.83 ;
      RECT  436.0025 192.55 436.4775 192.83 ;
      RECT  437.1775 192.55 437.6525 192.83 ;
      RECT  438.3525 192.55 438.8275 192.83 ;
      RECT  439.5275 192.55 440.0025 192.83 ;
      RECT  440.7025 192.55 441.1775 192.83 ;
      RECT  441.8775 192.55 442.3525 192.83 ;
      RECT  443.0525 192.55 443.5275 192.83 ;
      RECT  444.2275 192.55 444.7025 192.83 ;
      RECT  445.4025 192.55 445.8775 192.83 ;
      RECT  446.5775 192.55 447.0525 192.83 ;
      RECT  447.7525 192.55 448.2275 192.83 ;
      RECT  448.9275 192.55 449.4025 192.83 ;
      RECT  450.1025 192.55 450.5775 192.83 ;
      RECT  451.2775 192.55 451.7525 192.83 ;
      RECT  452.4525 192.55 452.9275 192.83 ;
      RECT  453.6275 192.55 454.1025 192.83 ;
      RECT  454.8025 192.55 455.2775 192.83 ;
      RECT  455.9775 192.55 456.4525 192.83 ;
      RECT  457.1525 192.55 457.6275 192.83 ;
      RECT  458.3275 192.55 458.8025 192.83 ;
      RECT  459.5025 192.55 459.9775 192.83 ;
      RECT  460.6775 192.55 461.1525 192.83 ;
      RECT  461.8525 192.55 462.3275 192.83 ;
      RECT  463.0275 192.55 463.5025 192.83 ;
      RECT  464.2025 192.55 464.6775 192.83 ;
      RECT  465.3775 192.55 465.8525 192.83 ;
      RECT  466.5525 192.55 467.0275 192.83 ;
      RECT  467.7275 192.55 468.2025 192.83 ;
      RECT  468.9025 192.55 469.3775 192.83 ;
      RECT  470.0775 192.55 470.5525 192.83 ;
      RECT  471.2525 192.55 471.7275 192.83 ;
      RECT  472.4275 192.55 472.9025 192.83 ;
      RECT  473.6025 192.55 474.0775 192.83 ;
      RECT  474.7775 192.55 475.2525 192.83 ;
      RECT  475.9525 192.55 476.4275 192.83 ;
      RECT  477.1275 192.55 477.6025 192.83 ;
      RECT  478.3025 192.55 478.7775 192.83 ;
      RECT  479.4775 192.55 479.9525 192.83 ;
      RECT  480.6525 192.55 481.1275 192.83 ;
      RECT  481.8275 192.55 482.3025 192.83 ;
      RECT  483.0025 192.55 483.4775 192.83 ;
      RECT  484.1775 192.55 484.6525 192.83 ;
      RECT  485.3525 192.55 485.8275 192.83 ;
      RECT  486.5275 192.55 487.0025 192.83 ;
      RECT  487.7025 192.55 488.1775 192.83 ;
      RECT  488.8775 192.55 489.3525 192.83 ;
      RECT  490.0525 192.55 490.5275 192.83 ;
      RECT  491.2275 192.55 491.7025 192.83 ;
      RECT  492.4025 192.55 492.8775 192.83 ;
      RECT  493.5775 192.55 494.0525 192.83 ;
      RECT  494.7525 192.55 495.2275 192.83 ;
      RECT  495.9275 192.55 496.4025 192.83 ;
      RECT  497.1025 192.55 497.5775 192.83 ;
      RECT  498.2775 192.55 498.7525 192.83 ;
      RECT  499.4525 192.55 499.9275 192.83 ;
      RECT  500.6275 192.55 501.1025 192.83 ;
      RECT  501.8025 192.55 502.2775 192.83 ;
      RECT  502.9775 192.55 503.4525 192.83 ;
      RECT  504.1525 192.55 504.6275 192.83 ;
      RECT  505.3275 192.55 505.8025 192.83 ;
      RECT  506.5025 192.55 506.9775 192.83 ;
      RECT  507.6775 192.55 508.1525 192.83 ;
      RECT  508.8525 192.55 509.3275 192.83 ;
      RECT  510.0275 192.55 510.5025 192.83 ;
      RECT  511.2025 192.55 511.6775 192.83 ;
      RECT  512.3775 192.55 512.8525 192.83 ;
      RECT  513.5525 192.55 514.0275 192.83 ;
      RECT  514.7275 192.55 515.2025 192.83 ;
      RECT  515.9025 192.55 516.3775 192.83 ;
      RECT  517.0775 192.55 517.5525 192.83 ;
      RECT  518.2525 192.55 518.7275 192.83 ;
      RECT  519.4275 192.55 519.9025 192.83 ;
      RECT  520.6025 192.55 521.0775 192.83 ;
      RECT  521.7775 192.55 522.2525 192.83 ;
      RECT  522.9525 192.55 523.4275 192.83 ;
      RECT  524.1275 192.55 524.6025 192.83 ;
      RECT  525.3025 192.55 525.7775 192.83 ;
      RECT  526.4775 192.55 526.9525 192.83 ;
      RECT  527.6525 192.55 528.1275 192.83 ;
      RECT  528.8275 192.55 529.3025 192.83 ;
      RECT  530.0025 192.55 530.4775 192.83 ;
      RECT  531.1775 192.55 531.6525 192.83 ;
      RECT  532.3525 192.55 532.8275 192.83 ;
      RECT  533.5275 192.55 534.0025 192.83 ;
      RECT  534.7025 192.55 535.1775 192.83 ;
      RECT  535.8775 192.55 536.3525 192.83 ;
      RECT  537.0525 192.55 537.5275 192.83 ;
      RECT  538.2275 192.55 538.7025 192.83 ;
      RECT  539.4025 192.55 539.8775 192.83 ;
      RECT  540.5775 192.55 541.0525 192.83 ;
      RECT  541.7525 192.55 542.2275 192.83 ;
      RECT  542.9275 192.55 543.4025 192.83 ;
      RECT  544.1025 192.55 544.5775 192.83 ;
      RECT  545.2775 192.55 545.7525 192.83 ;
      RECT  546.4525 192.55 546.9275 192.83 ;
      RECT  547.6275 192.55 548.1025 192.83 ;
      RECT  548.8025 192.55 549.2775 192.83 ;
      RECT  549.9775 192.55 550.4525 192.83 ;
      RECT  551.1525 192.55 551.6275 192.83 ;
      RECT  552.3275 192.55 552.8025 192.83 ;
      RECT  553.5025 192.55 553.9775 192.83 ;
      RECT  554.6775 192.55 555.1525 192.83 ;
      RECT  555.8525 192.55 556.3275 192.83 ;
      RECT  557.0275 192.55 557.5025 192.83 ;
      RECT  558.2025 192.55 558.6775 192.83 ;
      RECT  559.3775 192.55 559.8525 192.83 ;
      RECT  560.5525 192.55 561.0275 192.83 ;
      RECT  561.7275 192.55 562.2025 192.83 ;
      RECT  562.9025 192.55 563.3775 192.83 ;
      RECT  564.0775 192.55 564.5525 192.83 ;
      RECT  565.2525 192.55 565.7275 192.83 ;
      RECT  566.4275 192.55 566.9025 192.83 ;
      RECT  567.6025 192.55 568.0775 192.83 ;
      RECT  568.7775 192.55 569.2525 192.83 ;
      RECT  569.9525 192.55 570.4275 192.83 ;
      RECT  571.1275 192.55 571.6025 192.83 ;
      RECT  572.3025 192.55 572.7775 192.83 ;
      RECT  573.4775 192.55 573.9525 192.83 ;
      RECT  574.6525 192.55 575.1275 192.83 ;
      RECT  575.8275 192.55 576.3025 192.83 ;
      RECT  577.0025 192.55 577.4775 192.83 ;
      RECT  578.1775 192.55 578.6525 192.83 ;
      RECT  579.3525 192.55 579.8275 192.83 ;
      RECT  580.5275 192.55 581.0025 192.83 ;
      RECT  581.7025 192.55 582.1775 192.83 ;
      RECT  582.8775 192.55 583.3525 192.83 ;
      RECT  584.0525 192.55 584.5275 192.83 ;
      RECT  585.2275 192.55 585.7025 192.83 ;
      RECT  586.4025 192.55 586.8775 192.83 ;
      RECT  587.5775 192.55 588.0525 192.83 ;
      RECT  588.7525 192.55 589.2275 192.83 ;
      RECT  589.9275 192.55 590.4025 192.83 ;
      RECT  591.1025 192.55 591.5775 192.83 ;
      RECT  592.2775 192.55 592.7525 192.83 ;
      RECT  593.4525 192.55 593.9275 192.83 ;
      RECT  594.6275 192.55 595.1025 192.83 ;
      RECT  595.8025 192.55 596.2775 192.83 ;
      RECT  596.9775 192.55 597.4525 192.83 ;
      RECT  598.1525 192.55 598.6275 192.83 ;
      RECT  599.3275 192.55 599.8025 192.83 ;
      RECT  600.5025 192.55 600.9775 192.83 ;
      RECT  601.6775 192.55 602.1525 192.83 ;
      RECT  602.8525 192.55 603.3275 192.83 ;
      RECT  604.0275 192.55 604.5025 192.83 ;
      RECT  605.2025 192.55 605.6775 192.83 ;
      RECT  606.3775 192.55 606.8525 192.83 ;
      RECT  607.5525 192.55 608.0275 192.83 ;
      RECT  608.7275 192.55 609.2025 192.83 ;
      RECT  609.9025 192.55 610.3775 192.83 ;
      RECT  611.0775 192.55 611.5525 192.83 ;
      RECT  612.2525 192.55 612.7275 192.83 ;
      RECT  613.4275 192.55 613.9025 192.83 ;
      RECT  614.6025 192.55 615.0775 192.83 ;
      RECT  615.7775 192.55 616.2525 192.83 ;
      RECT  616.9525 192.55 617.4275 192.83 ;
      RECT  618.1275 192.55 618.6025 192.83 ;
      RECT  619.3025 192.55 619.7775 192.83 ;
      RECT  620.4775 192.55 620.9525 192.83 ;
      RECT  621.6525 192.55 622.1275 192.83 ;
      RECT  622.8275 192.55 623.3025 192.83 ;
      RECT  624.0025 192.55 624.4775 192.83 ;
      RECT  625.1775 192.55 625.6525 192.83 ;
      RECT  626.3525 192.55 626.8275 192.83 ;
      RECT  627.5275 192.55 628.0025 192.83 ;
      RECT  628.7025 192.55 629.1775 192.83 ;
      RECT  629.8775 192.55 630.3525 192.83 ;
      RECT  631.0525 192.55 631.5275 192.83 ;
      RECT  632.2275 192.55 632.7025 192.83 ;
      RECT  633.4025 192.55 633.8775 192.83 ;
      RECT  634.5775 192.55 635.0525 192.83 ;
      RECT  635.7525 192.55 636.2275 192.83 ;
      RECT  636.9275 192.55 637.4025 192.83 ;
      RECT  638.1025 192.55 638.5775 192.83 ;
      RECT  639.2775 192.55 639.7525 192.83 ;
      RECT  640.4525 192.55 640.9275 192.83 ;
      RECT  641.6275 192.55 642.1025 192.83 ;
      RECT  642.8025 192.55 643.2775 192.83 ;
      RECT  643.9775 192.55 644.4525 192.83 ;
      RECT  645.1525 192.55 645.6275 192.83 ;
      RECT  646.3275 192.55 646.8025 192.83 ;
      RECT  647.5025 192.55 647.9775 192.83 ;
      RECT  648.6775 192.55 649.1525 192.83 ;
      RECT  649.8525 192.55 650.3275 192.83 ;
      RECT  651.0275 192.55 651.5025 192.83 ;
      RECT  652.2025 192.55 652.6775 192.83 ;
      RECT  653.3775 192.55 653.8525 192.83 ;
      RECT  654.5525 192.55 655.0275 192.83 ;
      RECT  655.7275 192.55 656.2025 192.83 ;
      RECT  656.9025 192.55 657.3775 192.83 ;
      RECT  658.0775 192.55 658.5525 192.83 ;
      RECT  659.2525 192.55 659.7275 192.83 ;
      RECT  660.4275 192.55 660.9025 192.83 ;
      RECT  661.6025 192.55 662.0775 192.83 ;
      RECT  662.7775 192.55 663.2525 192.83 ;
      RECT  663.9525 192.55 664.4275 192.83 ;
      RECT  665.1275 192.55 665.6025 192.83 ;
      RECT  666.3025 192.55 666.7775 192.83 ;
      RECT  667.4775 192.55 667.9525 192.83 ;
      RECT  668.6525 192.55 669.1275 192.83 ;
      RECT  669.8275 192.55 670.3025 192.83 ;
      RECT  671.0025 192.55 671.4775 192.83 ;
      RECT  672.1775 192.55 672.6525 192.83 ;
      RECT  673.3525 192.55 673.8275 192.83 ;
      RECT  674.5275 192.55 675.0025 192.83 ;
      RECT  675.7025 192.55 676.1775 192.83 ;
      RECT  676.8775 192.55 677.3525 192.83 ;
      RECT  678.0525 192.55 678.5275 192.83 ;
      RECT  679.2275 192.55 679.7025 192.83 ;
      RECT  680.4025 192.55 680.8775 192.83 ;
      RECT  681.5775 192.55 682.0525 192.83 ;
      RECT  682.7525 192.55 683.2275 192.83 ;
      RECT  683.9275 192.55 684.4025 192.83 ;
      RECT  685.1025 192.55 685.5775 192.83 ;
      RECT  686.2775 192.55 686.7525 192.83 ;
      RECT  687.4525 192.55 687.9275 192.83 ;
      RECT  688.6275 192.55 689.1025 192.83 ;
      RECT  689.8025 192.55 690.2775 192.83 ;
      RECT  690.9775 192.55 691.4525 192.83 ;
      RECT  692.1525 192.55 692.6275 192.83 ;
      RECT  693.3275 192.55 693.8025 192.83 ;
      RECT  694.5025 192.55 694.9775 192.83 ;
      RECT  695.6775 192.55 696.1525 192.83 ;
      RECT  696.8525 192.55 697.3275 192.83 ;
      RECT  698.0275 192.55 698.5025 192.83 ;
      RECT  699.2025 192.55 699.6775 192.83 ;
      RECT  700.3775 192.55 700.8525 192.83 ;
      RECT  701.5525 192.55 702.0275 192.83 ;
      RECT  702.7275 192.55 703.2025 192.83 ;
      RECT  703.9025 192.55 704.3775 192.83 ;
      RECT  705.0775 192.55 705.5525 192.83 ;
      RECT  706.2525 192.55 706.7275 192.83 ;
      RECT  707.4275 192.55 707.9025 192.83 ;
      RECT  708.6025 192.55 709.0775 192.83 ;
      RECT  709.7775 192.55 710.2525 192.83 ;
      RECT  710.9525 192.55 711.4275 192.83 ;
      RECT  712.1275 192.55 712.6025 192.83 ;
      RECT  713.3025 192.55 713.7775 192.83 ;
      RECT  714.4775 192.55 714.9525 192.83 ;
      RECT  715.6525 192.55 716.1275 192.83 ;
      RECT  716.8275 192.55 717.3025 192.83 ;
      RECT  718.0025 192.55 718.4775 192.83 ;
      RECT  719.1775 192.55 719.6525 192.83 ;
      RECT  720.3525 192.55 720.8275 192.83 ;
      RECT  721.5275 192.55 722.0025 192.83 ;
      RECT  722.7025 192.55 723.1775 192.83 ;
      RECT  723.8775 192.55 724.3525 192.83 ;
      RECT  725.0525 192.55 725.5275 192.83 ;
      RECT  726.2275 192.55 726.7025 192.83 ;
      RECT  727.4025 192.55 727.8775 192.83 ;
      RECT  728.5775 192.55 729.0525 192.83 ;
      RECT  729.7525 192.55 730.2275 192.83 ;
      RECT  730.9275 192.55 731.4025 192.83 ;
      RECT  732.1025 192.55 732.5775 192.83 ;
      RECT  733.2775 192.55 733.7525 192.83 ;
      RECT  734.4525 192.55 734.9275 192.83 ;
      RECT  735.6275 192.55 736.1025 192.83 ;
      RECT  736.8025 192.55 737.2775 192.83 ;
      RECT  737.9775 192.55 738.4525 192.83 ;
      RECT  739.1525 192.55 739.6275 192.83 ;
      RECT  740.3275 192.55 740.8025 192.83 ;
      RECT  741.5025 192.55 741.9775 192.83 ;
      RECT  742.6775 192.55 743.1525 192.83 ;
      RECT  743.8525 192.55 744.3275 192.83 ;
      RECT  745.0275 192.55 745.5025 192.83 ;
      RECT  746.2025 192.55 746.6775 192.83 ;
      RECT  747.3775 192.55 747.8525 192.83 ;
      RECT  748.5525 192.55 749.0275 192.83 ;
      RECT  749.7275 192.55 750.2025 192.83 ;
      RECT  750.9025 192.55 751.3775 192.83 ;
      RECT  752.0775 192.55 752.5525 192.83 ;
      RECT  753.2525 192.55 753.7275 192.83 ;
      RECT  754.4275 192.55 754.9025 192.83 ;
      RECT  755.6025 192.55 756.0775 192.83 ;
      RECT  756.7775 192.55 757.2525 192.83 ;
      RECT  757.9525 192.55 758.4275 192.83 ;
      RECT  759.1275 192.55 759.6025 192.83 ;
      RECT  760.3025 192.55 760.7775 192.83 ;
      RECT  761.4775 192.55 761.9525 192.83 ;
      RECT  762.6525 192.55 763.1275 192.83 ;
      RECT  763.8275 192.55 764.3025 192.83 ;
      RECT  765.0025 192.55 765.4775 192.83 ;
      RECT  766.1775 192.55 766.6525 192.83 ;
      RECT  767.3525 192.55 767.8275 192.83 ;
      RECT  768.5275 192.55 769.0025 192.83 ;
      RECT  769.7025 192.55 770.1775 192.83 ;
      RECT  770.8775 192.55 771.3525 192.83 ;
      RECT  772.0525 192.55 772.5275 192.83 ;
      RECT  773.2275 192.55 773.7025 192.83 ;
      RECT  774.4025 192.55 774.8775 192.83 ;
      RECT  775.5775 192.55 776.0525 192.83 ;
      RECT  776.7525 192.55 777.2275 192.83 ;
      RECT  777.9275 192.55 778.4025 192.83 ;
      RECT  779.1025 192.55 779.5775 192.83 ;
      RECT  780.2775 192.55 780.7525 192.83 ;
      RECT  781.4525 192.55 781.9275 192.83 ;
      RECT  782.6275 192.55 783.1025 192.83 ;
      RECT  783.8025 192.55 784.2775 192.83 ;
      RECT  784.9775 192.55 785.4525 192.83 ;
      RECT  786.1525 192.55 786.6275 192.83 ;
      RECT  787.3275 192.55 787.8025 192.83 ;
      RECT  788.5025 192.55 788.9775 192.83 ;
      RECT  789.6775 192.55 790.1525 192.83 ;
      RECT  790.8525 192.55 791.3275 192.83 ;
      RECT  792.0275 192.55 792.5025 192.83 ;
      RECT  793.2025 192.55 793.6775 192.83 ;
      RECT  794.3775 192.55 794.8525 192.83 ;
      RECT  795.5525 192.55 796.0275 192.83 ;
      RECT  796.7275 192.55 797.2025 192.83 ;
      RECT  797.9025 192.55 798.3775 192.83 ;
      RECT  799.0775 192.55 799.5525 192.83 ;
      RECT  800.2525 192.55 800.7275 192.83 ;
      RECT  801.4275 192.55 801.9025 192.83 ;
      RECT  802.6025 192.55 803.0775 192.83 ;
      RECT  803.7775 192.55 804.2525 192.83 ;
      RECT  804.9525 192.55 805.4275 192.83 ;
      RECT  806.1275 192.55 806.6025 192.83 ;
      RECT  807.3025 192.55 807.7775 192.83 ;
      RECT  808.4775 192.55 808.9525 192.83 ;
      RECT  809.6525 192.55 810.1275 192.83 ;
      RECT  810.8275 192.55 811.3025 192.83 ;
      RECT  812.0025 192.55 812.4775 192.83 ;
      RECT  813.1775 192.55 813.6525 192.83 ;
      RECT  814.3525 192.55 814.8275 192.83 ;
      RECT  815.5275 192.55 816.0025 192.83 ;
      RECT  816.7025 192.55 817.1775 192.83 ;
      RECT  817.8775 192.55 818.3525 192.83 ;
      RECT  819.0525 192.55 819.5275 192.83 ;
      RECT  820.2275 192.55 820.7025 192.83 ;
      RECT  821.4025 192.55 821.8775 192.83 ;
      RECT  822.5775 192.55 823.0525 192.83 ;
      RECT  823.7525 192.55 824.2275 192.83 ;
      RECT  824.9275 192.55 825.4025 192.83 ;
      RECT  826.1025 192.55 826.5775 192.83 ;
      RECT  827.2775 192.55 827.7525 192.83 ;
      RECT  828.4525 192.55 828.9275 192.83 ;
      RECT  829.6275 192.55 830.1025 192.83 ;
      RECT  830.8025 192.55 831.2775 192.83 ;
      RECT  831.9775 192.55 832.4525 192.83 ;
      RECT  833.1525 192.55 833.6275 192.83 ;
      RECT  834.3275 192.55 834.8025 192.83 ;
      RECT  835.5025 192.55 835.9775 192.83 ;
      RECT  836.6775 192.55 837.1525 192.83 ;
      RECT  837.8525 192.55 838.3275 192.83 ;
      RECT  839.0275 192.55 839.5025 192.83 ;
      RECT  840.2025 192.55 840.6775 192.83 ;
      RECT  841.3775 192.55 841.8525 192.83 ;
      RECT  842.5525 192.55 843.0275 192.83 ;
      RECT  843.7275 192.55 844.2025 192.83 ;
      RECT  844.9025 192.55 845.3775 192.83 ;
      RECT  846.0775 192.55 846.5525 192.83 ;
      RECT  847.2525 192.55 847.7275 192.83 ;
      RECT  848.4275 192.55 848.9025 192.83 ;
      RECT  849.6025 192.55 891.065 192.83 ;
   END
END    sram_0rw1r1w_576_16_freepdk45
END    LIBRARY
