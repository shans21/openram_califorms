**************************************************
* OpenRAM generated memory.
* Words: 1024
* Data bits: 32
* Banks: 1
* Column mux: 8:1
* Trimmed: True
* LVS: False
**************************************************
* File: DFFPOSX1.pex.netlist
* Created: Wed Jan  2 18:36:24 2008
* Program "Calibre xRC"
* Version "v2007.2_34.24"
*
.subckt dff D Q clk vdd gnd
*
MM21 Q a_66_6# gnd gnd NMOS_VTG L=5e-08 W=5e-07
MM19 a_76_6# a_2_6# a_66_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM20 gnd Q a_76_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM18 a_66_6# clk a_61_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM17 a_61_6# a_34_4# gnd gnd NMOS_VTG L=5e-08 W=2.5e-07
MM10 gnd clk a_2_6# gnd NMOS_VTG L=5e-08 W=5e-07
MM16 a_34_4# a_22_6# gnd gnd NMOS_VTG L=5e-08 W=2.5e-07
MM15 gnd a_34_4# a_31_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM14 a_31_6# clk a_22_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM13 a_22_6# a_2_6# a_17_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM12 a_17_6# D gnd gnd NMOS_VTG L=5e-08 W=2.5e-07
MM11 Q a_66_6# vdd vdd PMOS_VTG L=5e-08 W=1e-06
MM9 vdd Q a_76_84# vdd PMOS_VTG L=5e-08 W=2.5e-07
MM8 a_76_84# clk a_66_6# vdd PMOS_VTG L=5e-08 W=2.5e-07
MM7 a_66_6# a_2_6# a_61_74# vdd PMOS_VTG L=5e-08 W=5e-07
MM6 a_61_74# a_34_4# vdd vdd PMOS_VTG L=5e-08 W=5e-07
MM0 vdd clk a_2_6# vdd PMOS_VTG L=5e-08 W=1e-06
MM5 a_34_4# a_22_6# vdd vdd PMOS_VTG L=5e-08 W=5e-07
MM4 vdd a_34_4# a_31_74# vdd PMOS_VTG L=5e-08 W=5e-07
MM3 a_31_74# a_2_6# a_22_6# vdd PMOS_VTG L=5e-08 W=5e-07
MM2 a_22_6# clk a_17_74# vdd PMOS_VTG L=5e-08 W=5e-07
MM1 a_17_74# D vdd vdd PMOS_VTG L=5e-08 W=5e-07
* c_9 a_66_6# 0 0.271997f
* c_20 clk 0 0.350944f
* c_27 Q 0 0.202617f
* c_32 a_76_84# 0 0.0210573f
* c_38 a_76_6# 0 0.0204911f
* c_45 a_34_4# 0 0.172306f
* c_55 a_2_6# 0 0.283119f
* c_59 a_22_6# 0 0.157312f
* c_64 D 0 0.0816386f
* c_73 gnd 0 0.254131f
* c_81 vdd 0 0.23624f
*
*.include "dff.pex.netlist.dff.pxi"
*
.ends
*
*

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_col_addr_dff
+ din_0 din_1 din_2 dout_0 dout_1 dout_2 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 3
Xdff_r0_c0
+ din_0 dout_0 clk vdd gnd
+ dff
Xdff_r0_c1
+ din_1 dout_1 clk vdd gnd
+ dff
Xdff_r0_c2
+ din_2 dout_2 clk vdd gnd
+ dff
.ENDS sram_1rw0r0w_32_1024_freepdk45_col_addr_dff

* spice ptx M{0} {1} nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p

* spice ptx M{0} {1} pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

* spice ptx M{0} {1} nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pnand2
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Mpnand2_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_nmos1 Z B net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand2_nmos2 net1 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pnand2

* spice ptx M{0} {1} nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p

* spice ptx M{0} {1} pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pinv
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pinv

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_and2_dec
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpand2_dec_nand
+ A B zb_int vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pnand2
Xpand2_dec_inv
+ zb_int Z vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv
.ENDS sram_1rw0r0w_32_1024_freepdk45_and2_dec

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_hierarchical_predecode2x4
+ in_0 in_1 out_0 out_1 out_2 out_3 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0
+ in_0 inbar_0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv
Xpre_inv_1
+ in_1 inbar_1 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv
XXpre2x4_and_0
+ inbar_0 inbar_1 out_0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and2_dec
XXpre2x4_and_1
+ in_0 inbar_1 out_1 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and2_dec
XXpre2x4_and_2
+ inbar_0 in_1 out_2 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and2_dec
XXpre2x4_and_3
+ in_0 in_1 out_3 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and2_dec
.ENDS sram_1rw0r0w_32_1024_freepdk45_hierarchical_predecode2x4

* spice ptx M{0} {1} nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pnand3
+ A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Mpnand3_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_pmos3 Z C vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_nmos1 Z C net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand3_nmos2 net1 B net2 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand3_nmos3 net2 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pnand3

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_and3_dec
+ A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpand3_dec_nand
+ A B C zb_int vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pnand3
Xpand3_dec_inv
+ zb_int Z vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv
.ENDS sram_1rw0r0w_32_1024_freepdk45_and3_dec

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_hierarchical_predecode3x8
+ in_0 in_1 in_2 out_0 out_1 out_2 out_3 out_4 out_5 out_6 out_7 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* OUTPUT: out_4 
* OUTPUT: out_5 
* OUTPUT: out_6 
* OUTPUT: out_7 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0
+ in_0 inbar_0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv
Xpre_inv_1
+ in_1 inbar_1 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv
Xpre_inv_2
+ in_2 inbar_2 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv
XXpre3x8_and_0
+ inbar_0 inbar_1 inbar_2 out_0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XXpre3x8_and_1
+ in_0 inbar_1 inbar_2 out_1 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XXpre3x8_and_2
+ inbar_0 in_1 inbar_2 out_2 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XXpre3x8_and_3
+ in_0 in_1 inbar_2 out_3 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XXpre3x8_and_4
+ inbar_0 inbar_1 in_2 out_4 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XXpre3x8_and_5
+ in_0 inbar_1 in_2 out_5 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XXpre3x8_and_6
+ inbar_0 in_1 in_2 out_6 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XXpre3x8_and_7
+ in_0 in_1 in_2 out_7 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
.ENDS sram_1rw0r0w_32_1024_freepdk45_hierarchical_predecode3x8

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_hierarchical_decoder
+ addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 addr_6 decode_0 decode_1
+ decode_2 decode_3 decode_4 decode_5 decode_6 decode_7 decode_8
+ decode_9 decode_10 decode_11 decode_12 decode_13 decode_14 decode_15
+ decode_16 decode_17 decode_18 decode_19 decode_20 decode_21 decode_22
+ decode_23 decode_24 decode_25 decode_26 decode_27 decode_28 decode_29
+ decode_30 decode_31 decode_32 decode_33 decode_34 decode_35 decode_36
+ decode_37 decode_38 decode_39 decode_40 decode_41 decode_42 decode_43
+ decode_44 decode_45 decode_46 decode_47 decode_48 decode_49 decode_50
+ decode_51 decode_52 decode_53 decode_54 decode_55 decode_56 decode_57
+ decode_58 decode_59 decode_60 decode_61 decode_62 decode_63 decode_64
+ decode_65 decode_66 decode_67 decode_68 decode_69 decode_70 decode_71
+ decode_72 decode_73 decode_74 decode_75 decode_76 decode_77 decode_78
+ decode_79 decode_80 decode_81 decode_82 decode_83 decode_84 decode_85
+ decode_86 decode_87 decode_88 decode_89 decode_90 decode_91 decode_92
+ decode_93 decode_94 decode_95 decode_96 decode_97 decode_98 decode_99
+ decode_100 decode_101 decode_102 decode_103 decode_104 decode_105
+ decode_106 decode_107 decode_108 decode_109 decode_110 decode_111
+ decode_112 decode_113 decode_114 decode_115 decode_116 decode_117
+ decode_118 decode_119 decode_120 decode_121 decode_122 decode_123
+ decode_124 decode_125 decode_126 decode_127 vdd gnd
* INPUT : addr_0 
* INPUT : addr_1 
* INPUT : addr_2 
* INPUT : addr_3 
* INPUT : addr_4 
* INPUT : addr_5 
* INPUT : addr_6 
* OUTPUT: decode_0 
* OUTPUT: decode_1 
* OUTPUT: decode_2 
* OUTPUT: decode_3 
* OUTPUT: decode_4 
* OUTPUT: decode_5 
* OUTPUT: decode_6 
* OUTPUT: decode_7 
* OUTPUT: decode_8 
* OUTPUT: decode_9 
* OUTPUT: decode_10 
* OUTPUT: decode_11 
* OUTPUT: decode_12 
* OUTPUT: decode_13 
* OUTPUT: decode_14 
* OUTPUT: decode_15 
* OUTPUT: decode_16 
* OUTPUT: decode_17 
* OUTPUT: decode_18 
* OUTPUT: decode_19 
* OUTPUT: decode_20 
* OUTPUT: decode_21 
* OUTPUT: decode_22 
* OUTPUT: decode_23 
* OUTPUT: decode_24 
* OUTPUT: decode_25 
* OUTPUT: decode_26 
* OUTPUT: decode_27 
* OUTPUT: decode_28 
* OUTPUT: decode_29 
* OUTPUT: decode_30 
* OUTPUT: decode_31 
* OUTPUT: decode_32 
* OUTPUT: decode_33 
* OUTPUT: decode_34 
* OUTPUT: decode_35 
* OUTPUT: decode_36 
* OUTPUT: decode_37 
* OUTPUT: decode_38 
* OUTPUT: decode_39 
* OUTPUT: decode_40 
* OUTPUT: decode_41 
* OUTPUT: decode_42 
* OUTPUT: decode_43 
* OUTPUT: decode_44 
* OUTPUT: decode_45 
* OUTPUT: decode_46 
* OUTPUT: decode_47 
* OUTPUT: decode_48 
* OUTPUT: decode_49 
* OUTPUT: decode_50 
* OUTPUT: decode_51 
* OUTPUT: decode_52 
* OUTPUT: decode_53 
* OUTPUT: decode_54 
* OUTPUT: decode_55 
* OUTPUT: decode_56 
* OUTPUT: decode_57 
* OUTPUT: decode_58 
* OUTPUT: decode_59 
* OUTPUT: decode_60 
* OUTPUT: decode_61 
* OUTPUT: decode_62 
* OUTPUT: decode_63 
* OUTPUT: decode_64 
* OUTPUT: decode_65 
* OUTPUT: decode_66 
* OUTPUT: decode_67 
* OUTPUT: decode_68 
* OUTPUT: decode_69 
* OUTPUT: decode_70 
* OUTPUT: decode_71 
* OUTPUT: decode_72 
* OUTPUT: decode_73 
* OUTPUT: decode_74 
* OUTPUT: decode_75 
* OUTPUT: decode_76 
* OUTPUT: decode_77 
* OUTPUT: decode_78 
* OUTPUT: decode_79 
* OUTPUT: decode_80 
* OUTPUT: decode_81 
* OUTPUT: decode_82 
* OUTPUT: decode_83 
* OUTPUT: decode_84 
* OUTPUT: decode_85 
* OUTPUT: decode_86 
* OUTPUT: decode_87 
* OUTPUT: decode_88 
* OUTPUT: decode_89 
* OUTPUT: decode_90 
* OUTPUT: decode_91 
* OUTPUT: decode_92 
* OUTPUT: decode_93 
* OUTPUT: decode_94 
* OUTPUT: decode_95 
* OUTPUT: decode_96 
* OUTPUT: decode_97 
* OUTPUT: decode_98 
* OUTPUT: decode_99 
* OUTPUT: decode_100 
* OUTPUT: decode_101 
* OUTPUT: decode_102 
* OUTPUT: decode_103 
* OUTPUT: decode_104 
* OUTPUT: decode_105 
* OUTPUT: decode_106 
* OUTPUT: decode_107 
* OUTPUT: decode_108 
* OUTPUT: decode_109 
* OUTPUT: decode_110 
* OUTPUT: decode_111 
* OUTPUT: decode_112 
* OUTPUT: decode_113 
* OUTPUT: decode_114 
* OUTPUT: decode_115 
* OUTPUT: decode_116 
* OUTPUT: decode_117 
* OUTPUT: decode_118 
* OUTPUT: decode_119 
* OUTPUT: decode_120 
* OUTPUT: decode_121 
* OUTPUT: decode_122 
* OUTPUT: decode_123 
* OUTPUT: decode_124 
* OUTPUT: decode_125 
* OUTPUT: decode_126 
* OUTPUT: decode_127 
* POWER : vdd 
* GROUND: gnd 
Xpre_0
+ addr_0 addr_1 out_0 out_1 out_2 out_3 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_hierarchical_predecode2x4
Xpre_1
+ addr_2 addr_3 out_4 out_5 out_6 out_7 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_hierarchical_predecode2x4
Xpre3x8_0
+ addr_4 addr_5 addr_6 out_8 out_9 out_10 out_11 out_12 out_13 out_14
+ out_15 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_hierarchical_predecode3x8
XDEC_AND_0
+ out_0 out_4 out_8 decode_0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_16
+ out_0 out_4 out_9 decode_16 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_32
+ out_0 out_4 out_10 decode_32 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_48
+ out_0 out_4 out_11 decode_48 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_64
+ out_0 out_4 out_12 decode_64 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_80
+ out_0 out_4 out_13 decode_80 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_96
+ out_0 out_4 out_14 decode_96 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_112
+ out_0 out_4 out_15 decode_112 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_4
+ out_0 out_5 out_8 decode_4 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_20
+ out_0 out_5 out_9 decode_20 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_36
+ out_0 out_5 out_10 decode_36 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_52
+ out_0 out_5 out_11 decode_52 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_68
+ out_0 out_5 out_12 decode_68 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_84
+ out_0 out_5 out_13 decode_84 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_100
+ out_0 out_5 out_14 decode_100 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_116
+ out_0 out_5 out_15 decode_116 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_8
+ out_0 out_6 out_8 decode_8 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_24
+ out_0 out_6 out_9 decode_24 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_40
+ out_0 out_6 out_10 decode_40 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_56
+ out_0 out_6 out_11 decode_56 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_72
+ out_0 out_6 out_12 decode_72 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_88
+ out_0 out_6 out_13 decode_88 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_104
+ out_0 out_6 out_14 decode_104 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_120
+ out_0 out_6 out_15 decode_120 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_12
+ out_0 out_7 out_8 decode_12 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_28
+ out_0 out_7 out_9 decode_28 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_44
+ out_0 out_7 out_10 decode_44 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_60
+ out_0 out_7 out_11 decode_60 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_76
+ out_0 out_7 out_12 decode_76 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_92
+ out_0 out_7 out_13 decode_92 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_108
+ out_0 out_7 out_14 decode_108 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_124
+ out_0 out_7 out_15 decode_124 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_1
+ out_1 out_4 out_8 decode_1 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_17
+ out_1 out_4 out_9 decode_17 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_33
+ out_1 out_4 out_10 decode_33 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_49
+ out_1 out_4 out_11 decode_49 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_65
+ out_1 out_4 out_12 decode_65 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_81
+ out_1 out_4 out_13 decode_81 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_97
+ out_1 out_4 out_14 decode_97 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_113
+ out_1 out_4 out_15 decode_113 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_5
+ out_1 out_5 out_8 decode_5 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_21
+ out_1 out_5 out_9 decode_21 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_37
+ out_1 out_5 out_10 decode_37 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_53
+ out_1 out_5 out_11 decode_53 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_69
+ out_1 out_5 out_12 decode_69 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_85
+ out_1 out_5 out_13 decode_85 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_101
+ out_1 out_5 out_14 decode_101 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_117
+ out_1 out_5 out_15 decode_117 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_9
+ out_1 out_6 out_8 decode_9 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_25
+ out_1 out_6 out_9 decode_25 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_41
+ out_1 out_6 out_10 decode_41 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_57
+ out_1 out_6 out_11 decode_57 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_73
+ out_1 out_6 out_12 decode_73 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_89
+ out_1 out_6 out_13 decode_89 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_105
+ out_1 out_6 out_14 decode_105 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_121
+ out_1 out_6 out_15 decode_121 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_13
+ out_1 out_7 out_8 decode_13 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_29
+ out_1 out_7 out_9 decode_29 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_45
+ out_1 out_7 out_10 decode_45 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_61
+ out_1 out_7 out_11 decode_61 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_77
+ out_1 out_7 out_12 decode_77 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_93
+ out_1 out_7 out_13 decode_93 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_109
+ out_1 out_7 out_14 decode_109 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_125
+ out_1 out_7 out_15 decode_125 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_2
+ out_2 out_4 out_8 decode_2 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_18
+ out_2 out_4 out_9 decode_18 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_34
+ out_2 out_4 out_10 decode_34 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_50
+ out_2 out_4 out_11 decode_50 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_66
+ out_2 out_4 out_12 decode_66 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_82
+ out_2 out_4 out_13 decode_82 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_98
+ out_2 out_4 out_14 decode_98 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_114
+ out_2 out_4 out_15 decode_114 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_6
+ out_2 out_5 out_8 decode_6 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_22
+ out_2 out_5 out_9 decode_22 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_38
+ out_2 out_5 out_10 decode_38 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_54
+ out_2 out_5 out_11 decode_54 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_70
+ out_2 out_5 out_12 decode_70 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_86
+ out_2 out_5 out_13 decode_86 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_102
+ out_2 out_5 out_14 decode_102 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_118
+ out_2 out_5 out_15 decode_118 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_10
+ out_2 out_6 out_8 decode_10 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_26
+ out_2 out_6 out_9 decode_26 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_42
+ out_2 out_6 out_10 decode_42 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_58
+ out_2 out_6 out_11 decode_58 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_74
+ out_2 out_6 out_12 decode_74 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_90
+ out_2 out_6 out_13 decode_90 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_106
+ out_2 out_6 out_14 decode_106 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_122
+ out_2 out_6 out_15 decode_122 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_14
+ out_2 out_7 out_8 decode_14 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_30
+ out_2 out_7 out_9 decode_30 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_46
+ out_2 out_7 out_10 decode_46 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_62
+ out_2 out_7 out_11 decode_62 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_78
+ out_2 out_7 out_12 decode_78 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_94
+ out_2 out_7 out_13 decode_94 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_110
+ out_2 out_7 out_14 decode_110 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_126
+ out_2 out_7 out_15 decode_126 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_3
+ out_3 out_4 out_8 decode_3 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_19
+ out_3 out_4 out_9 decode_19 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_35
+ out_3 out_4 out_10 decode_35 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_51
+ out_3 out_4 out_11 decode_51 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_67
+ out_3 out_4 out_12 decode_67 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_83
+ out_3 out_4 out_13 decode_83 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_99
+ out_3 out_4 out_14 decode_99 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_115
+ out_3 out_4 out_15 decode_115 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_7
+ out_3 out_5 out_8 decode_7 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_23
+ out_3 out_5 out_9 decode_23 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_39
+ out_3 out_5 out_10 decode_39 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_55
+ out_3 out_5 out_11 decode_55 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_71
+ out_3 out_5 out_12 decode_71 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_87
+ out_3 out_5 out_13 decode_87 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_103
+ out_3 out_5 out_14 decode_103 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_119
+ out_3 out_5 out_15 decode_119 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_11
+ out_3 out_6 out_8 decode_11 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_27
+ out_3 out_6 out_9 decode_27 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_43
+ out_3 out_6 out_10 decode_43 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_59
+ out_3 out_6 out_11 decode_59 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_75
+ out_3 out_6 out_12 decode_75 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_91
+ out_3 out_6 out_13 decode_91 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_107
+ out_3 out_6 out_14 decode_107 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_123
+ out_3 out_6 out_15 decode_123 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_15
+ out_3 out_7 out_8 decode_15 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_31
+ out_3 out_7 out_9 decode_31 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_47
+ out_3 out_7 out_10 decode_47 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_63
+ out_3 out_7 out_11 decode_63 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_79
+ out_3 out_7 out_12 decode_79 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_95
+ out_3 out_7 out_13 decode_95 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_111
+ out_3 out_7 out_14 decode_111 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
XDEC_AND_127
+ out_3 out_7 out_15 decode_127 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and3_dec
.ENDS sram_1rw0r0w_32_1024_freepdk45_hierarchical_decoder

* spice ptx M{0} {1} nmos_vtg m=47 w=0.1225u l=0.05u pd=0.34u ps=0.34u as=0.02p ad=0.02p

* spice ptx M{0} {1} pmos_vtg m=47 w=0.3675u l=0.05u pd=0.83u ps=0.83u as=0.05p ad=0.05p

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pinv_0
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 64
Mpinv_pmos Z A vdd vdd pmos_vtg m=47 w=0.3675u l=0.05u pd=0.83u ps=0.83u as=0.05p ad=0.05p
Mpinv_nmos Z A gnd gnd nmos_vtg m=47 w=0.1225u l=0.05u pd=0.34u ps=0.34u as=0.02p ad=0.02p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pinv_0

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_and2_dec_0
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 64
Xpand2_dec_nand
+ A B zb_int vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pnand2
Xpand2_dec_inv
+ zb_int Z vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_0
.ENDS sram_1rw0r0w_32_1024_freepdk45_and2_dec_0

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_wordline_driver
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* cols: 256
Xwld_nand
+ A B zb_int vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pnand2
Xwl_driver
+ zb_int Z vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_0
.ENDS sram_1rw0r0w_32_1024_freepdk45_wordline_driver

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_wordline_driver_array
+ in_0 in_1 in_2 in_3 in_4 in_5 in_6 in_7 in_8 in_9 in_10 in_11 in_12
+ in_13 in_14 in_15 in_16 in_17 in_18 in_19 in_20 in_21 in_22 in_23
+ in_24 in_25 in_26 in_27 in_28 in_29 in_30 in_31 in_32 in_33 in_34
+ in_35 in_36 in_37 in_38 in_39 in_40 in_41 in_42 in_43 in_44 in_45
+ in_46 in_47 in_48 in_49 in_50 in_51 in_52 in_53 in_54 in_55 in_56
+ in_57 in_58 in_59 in_60 in_61 in_62 in_63 in_64 in_65 in_66 in_67
+ in_68 in_69 in_70 in_71 in_72 in_73 in_74 in_75 in_76 in_77 in_78
+ in_79 in_80 in_81 in_82 in_83 in_84 in_85 in_86 in_87 in_88 in_89
+ in_90 in_91 in_92 in_93 in_94 in_95 in_96 in_97 in_98 in_99 in_100
+ in_101 in_102 in_103 in_104 in_105 in_106 in_107 in_108 in_109 in_110
+ in_111 in_112 in_113 in_114 in_115 in_116 in_117 in_118 in_119 in_120
+ in_121 in_122 in_123 in_124 in_125 in_126 in_127 wl_0 wl_1 wl_2 wl_3
+ wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15
+ wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26
+ wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37
+ wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48
+ wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59
+ wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70
+ wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81
+ wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92
+ wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103
+ wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113
+ wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123
+ wl_124 wl_125 wl_126 wl_127 en vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* INPUT : in_3 
* INPUT : in_4 
* INPUT : in_5 
* INPUT : in_6 
* INPUT : in_7 
* INPUT : in_8 
* INPUT : in_9 
* INPUT : in_10 
* INPUT : in_11 
* INPUT : in_12 
* INPUT : in_13 
* INPUT : in_14 
* INPUT : in_15 
* INPUT : in_16 
* INPUT : in_17 
* INPUT : in_18 
* INPUT : in_19 
* INPUT : in_20 
* INPUT : in_21 
* INPUT : in_22 
* INPUT : in_23 
* INPUT : in_24 
* INPUT : in_25 
* INPUT : in_26 
* INPUT : in_27 
* INPUT : in_28 
* INPUT : in_29 
* INPUT : in_30 
* INPUT : in_31 
* INPUT : in_32 
* INPUT : in_33 
* INPUT : in_34 
* INPUT : in_35 
* INPUT : in_36 
* INPUT : in_37 
* INPUT : in_38 
* INPUT : in_39 
* INPUT : in_40 
* INPUT : in_41 
* INPUT : in_42 
* INPUT : in_43 
* INPUT : in_44 
* INPUT : in_45 
* INPUT : in_46 
* INPUT : in_47 
* INPUT : in_48 
* INPUT : in_49 
* INPUT : in_50 
* INPUT : in_51 
* INPUT : in_52 
* INPUT : in_53 
* INPUT : in_54 
* INPUT : in_55 
* INPUT : in_56 
* INPUT : in_57 
* INPUT : in_58 
* INPUT : in_59 
* INPUT : in_60 
* INPUT : in_61 
* INPUT : in_62 
* INPUT : in_63 
* INPUT : in_64 
* INPUT : in_65 
* INPUT : in_66 
* INPUT : in_67 
* INPUT : in_68 
* INPUT : in_69 
* INPUT : in_70 
* INPUT : in_71 
* INPUT : in_72 
* INPUT : in_73 
* INPUT : in_74 
* INPUT : in_75 
* INPUT : in_76 
* INPUT : in_77 
* INPUT : in_78 
* INPUT : in_79 
* INPUT : in_80 
* INPUT : in_81 
* INPUT : in_82 
* INPUT : in_83 
* INPUT : in_84 
* INPUT : in_85 
* INPUT : in_86 
* INPUT : in_87 
* INPUT : in_88 
* INPUT : in_89 
* INPUT : in_90 
* INPUT : in_91 
* INPUT : in_92 
* INPUT : in_93 
* INPUT : in_94 
* INPUT : in_95 
* INPUT : in_96 
* INPUT : in_97 
* INPUT : in_98 
* INPUT : in_99 
* INPUT : in_100 
* INPUT : in_101 
* INPUT : in_102 
* INPUT : in_103 
* INPUT : in_104 
* INPUT : in_105 
* INPUT : in_106 
* INPUT : in_107 
* INPUT : in_108 
* INPUT : in_109 
* INPUT : in_110 
* INPUT : in_111 
* INPUT : in_112 
* INPUT : in_113 
* INPUT : in_114 
* INPUT : in_115 
* INPUT : in_116 
* INPUT : in_117 
* INPUT : in_118 
* INPUT : in_119 
* INPUT : in_120 
* INPUT : in_121 
* INPUT : in_122 
* INPUT : in_123 
* INPUT : in_124 
* INPUT : in_125 
* INPUT : in_126 
* INPUT : in_127 
* OUTPUT: wl_0 
* OUTPUT: wl_1 
* OUTPUT: wl_2 
* OUTPUT: wl_3 
* OUTPUT: wl_4 
* OUTPUT: wl_5 
* OUTPUT: wl_6 
* OUTPUT: wl_7 
* OUTPUT: wl_8 
* OUTPUT: wl_9 
* OUTPUT: wl_10 
* OUTPUT: wl_11 
* OUTPUT: wl_12 
* OUTPUT: wl_13 
* OUTPUT: wl_14 
* OUTPUT: wl_15 
* OUTPUT: wl_16 
* OUTPUT: wl_17 
* OUTPUT: wl_18 
* OUTPUT: wl_19 
* OUTPUT: wl_20 
* OUTPUT: wl_21 
* OUTPUT: wl_22 
* OUTPUT: wl_23 
* OUTPUT: wl_24 
* OUTPUT: wl_25 
* OUTPUT: wl_26 
* OUTPUT: wl_27 
* OUTPUT: wl_28 
* OUTPUT: wl_29 
* OUTPUT: wl_30 
* OUTPUT: wl_31 
* OUTPUT: wl_32 
* OUTPUT: wl_33 
* OUTPUT: wl_34 
* OUTPUT: wl_35 
* OUTPUT: wl_36 
* OUTPUT: wl_37 
* OUTPUT: wl_38 
* OUTPUT: wl_39 
* OUTPUT: wl_40 
* OUTPUT: wl_41 
* OUTPUT: wl_42 
* OUTPUT: wl_43 
* OUTPUT: wl_44 
* OUTPUT: wl_45 
* OUTPUT: wl_46 
* OUTPUT: wl_47 
* OUTPUT: wl_48 
* OUTPUT: wl_49 
* OUTPUT: wl_50 
* OUTPUT: wl_51 
* OUTPUT: wl_52 
* OUTPUT: wl_53 
* OUTPUT: wl_54 
* OUTPUT: wl_55 
* OUTPUT: wl_56 
* OUTPUT: wl_57 
* OUTPUT: wl_58 
* OUTPUT: wl_59 
* OUTPUT: wl_60 
* OUTPUT: wl_61 
* OUTPUT: wl_62 
* OUTPUT: wl_63 
* OUTPUT: wl_64 
* OUTPUT: wl_65 
* OUTPUT: wl_66 
* OUTPUT: wl_67 
* OUTPUT: wl_68 
* OUTPUT: wl_69 
* OUTPUT: wl_70 
* OUTPUT: wl_71 
* OUTPUT: wl_72 
* OUTPUT: wl_73 
* OUTPUT: wl_74 
* OUTPUT: wl_75 
* OUTPUT: wl_76 
* OUTPUT: wl_77 
* OUTPUT: wl_78 
* OUTPUT: wl_79 
* OUTPUT: wl_80 
* OUTPUT: wl_81 
* OUTPUT: wl_82 
* OUTPUT: wl_83 
* OUTPUT: wl_84 
* OUTPUT: wl_85 
* OUTPUT: wl_86 
* OUTPUT: wl_87 
* OUTPUT: wl_88 
* OUTPUT: wl_89 
* OUTPUT: wl_90 
* OUTPUT: wl_91 
* OUTPUT: wl_92 
* OUTPUT: wl_93 
* OUTPUT: wl_94 
* OUTPUT: wl_95 
* OUTPUT: wl_96 
* OUTPUT: wl_97 
* OUTPUT: wl_98 
* OUTPUT: wl_99 
* OUTPUT: wl_100 
* OUTPUT: wl_101 
* OUTPUT: wl_102 
* OUTPUT: wl_103 
* OUTPUT: wl_104 
* OUTPUT: wl_105 
* OUTPUT: wl_106 
* OUTPUT: wl_107 
* OUTPUT: wl_108 
* OUTPUT: wl_109 
* OUTPUT: wl_110 
* OUTPUT: wl_111 
* OUTPUT: wl_112 
* OUTPUT: wl_113 
* OUTPUT: wl_114 
* OUTPUT: wl_115 
* OUTPUT: wl_116 
* OUTPUT: wl_117 
* OUTPUT: wl_118 
* OUTPUT: wl_119 
* OUTPUT: wl_120 
* OUTPUT: wl_121 
* OUTPUT: wl_122 
* OUTPUT: wl_123 
* OUTPUT: wl_124 
* OUTPUT: wl_125 
* OUTPUT: wl_126 
* OUTPUT: wl_127 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* rows: 128 cols: 256
Xwl_driver_and0
+ in_0 en wl_0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and1
+ in_1 en wl_1 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and2
+ in_2 en wl_2 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and3
+ in_3 en wl_3 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and4
+ in_4 en wl_4 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and5
+ in_5 en wl_5 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and6
+ in_6 en wl_6 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and7
+ in_7 en wl_7 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and8
+ in_8 en wl_8 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and9
+ in_9 en wl_9 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and10
+ in_10 en wl_10 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and11
+ in_11 en wl_11 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and12
+ in_12 en wl_12 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and13
+ in_13 en wl_13 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and14
+ in_14 en wl_14 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and15
+ in_15 en wl_15 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and16
+ in_16 en wl_16 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and17
+ in_17 en wl_17 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and18
+ in_18 en wl_18 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and19
+ in_19 en wl_19 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and20
+ in_20 en wl_20 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and21
+ in_21 en wl_21 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and22
+ in_22 en wl_22 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and23
+ in_23 en wl_23 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and24
+ in_24 en wl_24 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and25
+ in_25 en wl_25 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and26
+ in_26 en wl_26 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and27
+ in_27 en wl_27 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and28
+ in_28 en wl_28 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and29
+ in_29 en wl_29 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and30
+ in_30 en wl_30 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and31
+ in_31 en wl_31 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and32
+ in_32 en wl_32 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and33
+ in_33 en wl_33 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and34
+ in_34 en wl_34 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and35
+ in_35 en wl_35 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and36
+ in_36 en wl_36 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and37
+ in_37 en wl_37 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and38
+ in_38 en wl_38 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and39
+ in_39 en wl_39 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and40
+ in_40 en wl_40 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and41
+ in_41 en wl_41 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and42
+ in_42 en wl_42 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and43
+ in_43 en wl_43 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and44
+ in_44 en wl_44 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and45
+ in_45 en wl_45 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and46
+ in_46 en wl_46 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and47
+ in_47 en wl_47 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and48
+ in_48 en wl_48 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and49
+ in_49 en wl_49 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and50
+ in_50 en wl_50 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and51
+ in_51 en wl_51 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and52
+ in_52 en wl_52 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and53
+ in_53 en wl_53 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and54
+ in_54 en wl_54 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and55
+ in_55 en wl_55 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and56
+ in_56 en wl_56 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and57
+ in_57 en wl_57 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and58
+ in_58 en wl_58 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and59
+ in_59 en wl_59 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and60
+ in_60 en wl_60 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and61
+ in_61 en wl_61 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and62
+ in_62 en wl_62 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and63
+ in_63 en wl_63 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and64
+ in_64 en wl_64 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and65
+ in_65 en wl_65 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and66
+ in_66 en wl_66 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and67
+ in_67 en wl_67 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and68
+ in_68 en wl_68 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and69
+ in_69 en wl_69 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and70
+ in_70 en wl_70 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and71
+ in_71 en wl_71 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and72
+ in_72 en wl_72 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and73
+ in_73 en wl_73 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and74
+ in_74 en wl_74 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and75
+ in_75 en wl_75 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and76
+ in_76 en wl_76 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and77
+ in_77 en wl_77 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and78
+ in_78 en wl_78 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and79
+ in_79 en wl_79 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and80
+ in_80 en wl_80 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and81
+ in_81 en wl_81 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and82
+ in_82 en wl_82 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and83
+ in_83 en wl_83 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and84
+ in_84 en wl_84 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and85
+ in_85 en wl_85 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and86
+ in_86 en wl_86 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and87
+ in_87 en wl_87 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and88
+ in_88 en wl_88 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and89
+ in_89 en wl_89 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and90
+ in_90 en wl_90 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and91
+ in_91 en wl_91 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and92
+ in_92 en wl_92 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and93
+ in_93 en wl_93 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and94
+ in_94 en wl_94 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and95
+ in_95 en wl_95 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and96
+ in_96 en wl_96 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and97
+ in_97 en wl_97 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and98
+ in_98 en wl_98 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and99
+ in_99 en wl_99 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and100
+ in_100 en wl_100 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and101
+ in_101 en wl_101 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and102
+ in_102 en wl_102 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and103
+ in_103 en wl_103 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and104
+ in_104 en wl_104 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and105
+ in_105 en wl_105 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and106
+ in_106 en wl_106 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and107
+ in_107 en wl_107 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and108
+ in_108 en wl_108 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and109
+ in_109 en wl_109 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and110
+ in_110 en wl_110 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and111
+ in_111 en wl_111 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and112
+ in_112 en wl_112 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and113
+ in_113 en wl_113 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and114
+ in_114 en wl_114 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and115
+ in_115 en wl_115 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and116
+ in_116 en wl_116 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and117
+ in_117 en wl_117 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and118
+ in_118 en wl_118 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and119
+ in_119 en wl_119 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and120
+ in_120 en wl_120 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and121
+ in_121 en wl_121 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and122
+ in_122 en wl_122 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and123
+ in_123 en wl_123 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and124
+ in_124 en wl_124 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and125
+ in_125 en wl_125 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and126
+ in_126 en wl_126 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
Xwl_driver_and127
+ in_127 en wl_127 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver
.ENDS sram_1rw0r0w_32_1024_freepdk45_wordline_driver_array

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_port_address
+ addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 addr_6 wl_en wl_0 wl_1 wl_2
+ wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15
+ wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26
+ wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37
+ wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48
+ wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59
+ wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70
+ wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81
+ wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92
+ wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103
+ wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113
+ wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123
+ wl_124 wl_125 wl_126 wl_127 rbl_wl vdd gnd
* INPUT : addr_0 
* INPUT : addr_1 
* INPUT : addr_2 
* INPUT : addr_3 
* INPUT : addr_4 
* INPUT : addr_5 
* INPUT : addr_6 
* INPUT : wl_en 
* OUTPUT: wl_0 
* OUTPUT: wl_1 
* OUTPUT: wl_2 
* OUTPUT: wl_3 
* OUTPUT: wl_4 
* OUTPUT: wl_5 
* OUTPUT: wl_6 
* OUTPUT: wl_7 
* OUTPUT: wl_8 
* OUTPUT: wl_9 
* OUTPUT: wl_10 
* OUTPUT: wl_11 
* OUTPUT: wl_12 
* OUTPUT: wl_13 
* OUTPUT: wl_14 
* OUTPUT: wl_15 
* OUTPUT: wl_16 
* OUTPUT: wl_17 
* OUTPUT: wl_18 
* OUTPUT: wl_19 
* OUTPUT: wl_20 
* OUTPUT: wl_21 
* OUTPUT: wl_22 
* OUTPUT: wl_23 
* OUTPUT: wl_24 
* OUTPUT: wl_25 
* OUTPUT: wl_26 
* OUTPUT: wl_27 
* OUTPUT: wl_28 
* OUTPUT: wl_29 
* OUTPUT: wl_30 
* OUTPUT: wl_31 
* OUTPUT: wl_32 
* OUTPUT: wl_33 
* OUTPUT: wl_34 
* OUTPUT: wl_35 
* OUTPUT: wl_36 
* OUTPUT: wl_37 
* OUTPUT: wl_38 
* OUTPUT: wl_39 
* OUTPUT: wl_40 
* OUTPUT: wl_41 
* OUTPUT: wl_42 
* OUTPUT: wl_43 
* OUTPUT: wl_44 
* OUTPUT: wl_45 
* OUTPUT: wl_46 
* OUTPUT: wl_47 
* OUTPUT: wl_48 
* OUTPUT: wl_49 
* OUTPUT: wl_50 
* OUTPUT: wl_51 
* OUTPUT: wl_52 
* OUTPUT: wl_53 
* OUTPUT: wl_54 
* OUTPUT: wl_55 
* OUTPUT: wl_56 
* OUTPUT: wl_57 
* OUTPUT: wl_58 
* OUTPUT: wl_59 
* OUTPUT: wl_60 
* OUTPUT: wl_61 
* OUTPUT: wl_62 
* OUTPUT: wl_63 
* OUTPUT: wl_64 
* OUTPUT: wl_65 
* OUTPUT: wl_66 
* OUTPUT: wl_67 
* OUTPUT: wl_68 
* OUTPUT: wl_69 
* OUTPUT: wl_70 
* OUTPUT: wl_71 
* OUTPUT: wl_72 
* OUTPUT: wl_73 
* OUTPUT: wl_74 
* OUTPUT: wl_75 
* OUTPUT: wl_76 
* OUTPUT: wl_77 
* OUTPUT: wl_78 
* OUTPUT: wl_79 
* OUTPUT: wl_80 
* OUTPUT: wl_81 
* OUTPUT: wl_82 
* OUTPUT: wl_83 
* OUTPUT: wl_84 
* OUTPUT: wl_85 
* OUTPUT: wl_86 
* OUTPUT: wl_87 
* OUTPUT: wl_88 
* OUTPUT: wl_89 
* OUTPUT: wl_90 
* OUTPUT: wl_91 
* OUTPUT: wl_92 
* OUTPUT: wl_93 
* OUTPUT: wl_94 
* OUTPUT: wl_95 
* OUTPUT: wl_96 
* OUTPUT: wl_97 
* OUTPUT: wl_98 
* OUTPUT: wl_99 
* OUTPUT: wl_100 
* OUTPUT: wl_101 
* OUTPUT: wl_102 
* OUTPUT: wl_103 
* OUTPUT: wl_104 
* OUTPUT: wl_105 
* OUTPUT: wl_106 
* OUTPUT: wl_107 
* OUTPUT: wl_108 
* OUTPUT: wl_109 
* OUTPUT: wl_110 
* OUTPUT: wl_111 
* OUTPUT: wl_112 
* OUTPUT: wl_113 
* OUTPUT: wl_114 
* OUTPUT: wl_115 
* OUTPUT: wl_116 
* OUTPUT: wl_117 
* OUTPUT: wl_118 
* OUTPUT: wl_119 
* OUTPUT: wl_120 
* OUTPUT: wl_121 
* OUTPUT: wl_122 
* OUTPUT: wl_123 
* OUTPUT: wl_124 
* OUTPUT: wl_125 
* OUTPUT: wl_126 
* OUTPUT: wl_127 
* OUTPUT: rbl_wl 
* POWER : vdd 
* GROUND: gnd 
Xrow_decoder
+ addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 addr_6 dec_out_0 dec_out_1
+ dec_out_2 dec_out_3 dec_out_4 dec_out_5 dec_out_6 dec_out_7 dec_out_8
+ dec_out_9 dec_out_10 dec_out_11 dec_out_12 dec_out_13 dec_out_14
+ dec_out_15 dec_out_16 dec_out_17 dec_out_18 dec_out_19 dec_out_20
+ dec_out_21 dec_out_22 dec_out_23 dec_out_24 dec_out_25 dec_out_26
+ dec_out_27 dec_out_28 dec_out_29 dec_out_30 dec_out_31 dec_out_32
+ dec_out_33 dec_out_34 dec_out_35 dec_out_36 dec_out_37 dec_out_38
+ dec_out_39 dec_out_40 dec_out_41 dec_out_42 dec_out_43 dec_out_44
+ dec_out_45 dec_out_46 dec_out_47 dec_out_48 dec_out_49 dec_out_50
+ dec_out_51 dec_out_52 dec_out_53 dec_out_54 dec_out_55 dec_out_56
+ dec_out_57 dec_out_58 dec_out_59 dec_out_60 dec_out_61 dec_out_62
+ dec_out_63 dec_out_64 dec_out_65 dec_out_66 dec_out_67 dec_out_68
+ dec_out_69 dec_out_70 dec_out_71 dec_out_72 dec_out_73 dec_out_74
+ dec_out_75 dec_out_76 dec_out_77 dec_out_78 dec_out_79 dec_out_80
+ dec_out_81 dec_out_82 dec_out_83 dec_out_84 dec_out_85 dec_out_86
+ dec_out_87 dec_out_88 dec_out_89 dec_out_90 dec_out_91 dec_out_92
+ dec_out_93 dec_out_94 dec_out_95 dec_out_96 dec_out_97 dec_out_98
+ dec_out_99 dec_out_100 dec_out_101 dec_out_102 dec_out_103 dec_out_104
+ dec_out_105 dec_out_106 dec_out_107 dec_out_108 dec_out_109
+ dec_out_110 dec_out_111 dec_out_112 dec_out_113 dec_out_114
+ dec_out_115 dec_out_116 dec_out_117 dec_out_118 dec_out_119
+ dec_out_120 dec_out_121 dec_out_122 dec_out_123 dec_out_124
+ dec_out_125 dec_out_126 dec_out_127 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_hierarchical_decoder
Xwordline_driver
+ dec_out_0 dec_out_1 dec_out_2 dec_out_3 dec_out_4 dec_out_5 dec_out_6
+ dec_out_7 dec_out_8 dec_out_9 dec_out_10 dec_out_11 dec_out_12
+ dec_out_13 dec_out_14 dec_out_15 dec_out_16 dec_out_17 dec_out_18
+ dec_out_19 dec_out_20 dec_out_21 dec_out_22 dec_out_23 dec_out_24
+ dec_out_25 dec_out_26 dec_out_27 dec_out_28 dec_out_29 dec_out_30
+ dec_out_31 dec_out_32 dec_out_33 dec_out_34 dec_out_35 dec_out_36
+ dec_out_37 dec_out_38 dec_out_39 dec_out_40 dec_out_41 dec_out_42
+ dec_out_43 dec_out_44 dec_out_45 dec_out_46 dec_out_47 dec_out_48
+ dec_out_49 dec_out_50 dec_out_51 dec_out_52 dec_out_53 dec_out_54
+ dec_out_55 dec_out_56 dec_out_57 dec_out_58 dec_out_59 dec_out_60
+ dec_out_61 dec_out_62 dec_out_63 dec_out_64 dec_out_65 dec_out_66
+ dec_out_67 dec_out_68 dec_out_69 dec_out_70 dec_out_71 dec_out_72
+ dec_out_73 dec_out_74 dec_out_75 dec_out_76 dec_out_77 dec_out_78
+ dec_out_79 dec_out_80 dec_out_81 dec_out_82 dec_out_83 dec_out_84
+ dec_out_85 dec_out_86 dec_out_87 dec_out_88 dec_out_89 dec_out_90
+ dec_out_91 dec_out_92 dec_out_93 dec_out_94 dec_out_95 dec_out_96
+ dec_out_97 dec_out_98 dec_out_99 dec_out_100 dec_out_101 dec_out_102
+ dec_out_103 dec_out_104 dec_out_105 dec_out_106 dec_out_107
+ dec_out_108 dec_out_109 dec_out_110 dec_out_111 dec_out_112
+ dec_out_113 dec_out_114 dec_out_115 dec_out_116 dec_out_117
+ dec_out_118 dec_out_119 dec_out_120 dec_out_121 dec_out_122
+ dec_out_123 dec_out_124 dec_out_125 dec_out_126 dec_out_127 wl_0 wl_1
+ wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14
+ wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25
+ wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36
+ wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47
+ wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58
+ wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69
+ wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80
+ wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91
+ wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102
+ wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112
+ wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122
+ wl_123 wl_124 wl_125 wl_126 wl_127 wl_en vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_wordline_driver_array
Xrbl_driver
+ wl_en vdd rbl_wl vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_and2_dec_0
.ENDS sram_1rw0r0w_32_1024_freepdk45_port_address

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pinv_2
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pinv_2

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pinv_1
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pinv_1

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pdriver
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1]
Xbuf_inv1
+ A Z vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_1
.ENDS sram_1rw0r0w_32_1024_freepdk45_pdriver

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pnand3_0
+ A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Mpnand3_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_pmos3 Z C vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_nmos1 Z C net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand3_nmos2 net1 B net2 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand3_nmos3 net2 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pnand3_0

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pand3
+ A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpand3_nand
+ A B C zb_int vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pnand3_0
Xpand3_inv
+ zb_int Z vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pdriver
.ENDS sram_1rw0r0w_32_1024_freepdk45_pand3

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_hierarchical_predecode3x8_0
+ in_0 in_1 in_2 out_0 out_1 out_2 out_3 out_4 out_5 out_6 out_7 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* OUTPUT: out_4 
* OUTPUT: out_5 
* OUTPUT: out_6 
* OUTPUT: out_7 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0
+ in_0 inbar_0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_2
Xpre_inv_1
+ in_1 inbar_1 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_2
Xpre_inv_2
+ in_2 inbar_2 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_2
XXpre3x8_and_0
+ inbar_0 inbar_1 inbar_2 out_0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pand3
XXpre3x8_and_1
+ in_0 inbar_1 inbar_2 out_1 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pand3
XXpre3x8_and_2
+ inbar_0 in_1 inbar_2 out_2 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pand3
XXpre3x8_and_3
+ in_0 in_1 inbar_2 out_3 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pand3
XXpre3x8_and_4
+ inbar_0 inbar_1 in_2 out_4 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pand3
XXpre3x8_and_5
+ in_0 inbar_1 in_2 out_5 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pand3
XXpre3x8_and_6
+ inbar_0 in_1 in_2 out_6 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pand3
XXpre3x8_and_7
+ in_0 in_1 in_2 out_7 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pand3
.ENDS sram_1rw0r0w_32_1024_freepdk45_hierarchical_predecode3x8_0

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_column_decoder
+ in_0 in_1 in_2 out_0 out_1 out_2 out_3 out_4 out_5 out_6 out_7 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* OUTPUT: out_4 
* OUTPUT: out_5 
* OUTPUT: out_6 
* OUTPUT: out_7 
* POWER : vdd 
* GROUND: gnd 
Xcolumn_decoder
+ in_0 in_1 in_2 out_0 out_1 out_2 out_3 out_4 out_5 out_6 out_7 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_hierarchical_predecode3x8_0
.ENDS sram_1rw0r0w_32_1024_freepdk45_column_decoder

.SUBCKT dummy_cell_1rw bl br wl vdd gnd
* Inverter 1
MM0 Q_bar Q gnd gnd NMOS_VTG W=205.00n L=50n
MM4 Q_bar Q vdd vdd PMOS_VTG W=90n L=50n

* Inverer 2
MM1 Q Q_bar gnd gnd NMOS_VTG W=205.00n L=50n
MM5 Q Q_bar vdd vdd PMOS_VTG W=90n L=50n

* Access transistors
MM3 bl_noconn wl Q gnd NMOS_VTG W=135.00n L=50n
MM2 br_noconn wl Q_bar gnd NMOS_VTG W=135.00n L=50n
.ENDS dummy_cell_1rw


.SUBCKT sram_1rw0r0w_32_1024_freepdk45_dummy_array_1
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65
+ bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69
+ bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73
+ bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77
+ bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81
+ bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85
+ bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89
+ bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93
+ bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97
+ bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101
+ bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105
+ br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108
+ bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112
+ br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115
+ bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119
+ br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122
+ bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126
+ br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 bl_0_129 br_0_129
+ bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132 br_0_132 bl_0_133
+ br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135 bl_0_136 br_0_136
+ bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139 br_0_139 bl_0_140
+ br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142 bl_0_143 br_0_143
+ bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146 br_0_146 bl_0_147
+ br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149 bl_0_150 br_0_150
+ bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153 br_0_153 bl_0_154
+ br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156 bl_0_157 br_0_157
+ bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160 br_0_160 bl_0_161
+ br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163 bl_0_164 br_0_164
+ bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167 br_0_167 bl_0_168
+ br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170 bl_0_171 br_0_171
+ bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174 br_0_174 bl_0_175
+ br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177 bl_0_178 br_0_178
+ bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181 br_0_181 bl_0_182
+ br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184 bl_0_185 br_0_185
+ bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188 br_0_188 bl_0_189
+ br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191 bl_0_192 br_0_192
+ bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195 br_0_195 bl_0_196
+ br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198 bl_0_199 br_0_199
+ bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202 br_0_202 bl_0_203
+ br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205 bl_0_206 br_0_206
+ bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209 br_0_209 bl_0_210
+ br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212 bl_0_213 br_0_213
+ bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216 br_0_216 bl_0_217
+ br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219 bl_0_220 br_0_220
+ bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223 br_0_223 bl_0_224
+ br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226 bl_0_227 br_0_227
+ bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230 br_0_230 bl_0_231
+ br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233 bl_0_234 br_0_234
+ bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237 br_0_237 bl_0_238
+ br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240 bl_0_241 br_0_241
+ bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244 br_0_244 bl_0_245
+ br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247 bl_0_248 br_0_248
+ bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251 br_0_251 bl_0_252
+ br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254 bl_0_255 br_0_255
+ bl_0_256 br_0_256 wl_0_0 vdd gnd
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INOUT : bl_0_64 
* INOUT : br_0_64 
* INOUT : bl_0_65 
* INOUT : br_0_65 
* INOUT : bl_0_66 
* INOUT : br_0_66 
* INOUT : bl_0_67 
* INOUT : br_0_67 
* INOUT : bl_0_68 
* INOUT : br_0_68 
* INOUT : bl_0_69 
* INOUT : br_0_69 
* INOUT : bl_0_70 
* INOUT : br_0_70 
* INOUT : bl_0_71 
* INOUT : br_0_71 
* INOUT : bl_0_72 
* INOUT : br_0_72 
* INOUT : bl_0_73 
* INOUT : br_0_73 
* INOUT : bl_0_74 
* INOUT : br_0_74 
* INOUT : bl_0_75 
* INOUT : br_0_75 
* INOUT : bl_0_76 
* INOUT : br_0_76 
* INOUT : bl_0_77 
* INOUT : br_0_77 
* INOUT : bl_0_78 
* INOUT : br_0_78 
* INOUT : bl_0_79 
* INOUT : br_0_79 
* INOUT : bl_0_80 
* INOUT : br_0_80 
* INOUT : bl_0_81 
* INOUT : br_0_81 
* INOUT : bl_0_82 
* INOUT : br_0_82 
* INOUT : bl_0_83 
* INOUT : br_0_83 
* INOUT : bl_0_84 
* INOUT : br_0_84 
* INOUT : bl_0_85 
* INOUT : br_0_85 
* INOUT : bl_0_86 
* INOUT : br_0_86 
* INOUT : bl_0_87 
* INOUT : br_0_87 
* INOUT : bl_0_88 
* INOUT : br_0_88 
* INOUT : bl_0_89 
* INOUT : br_0_89 
* INOUT : bl_0_90 
* INOUT : br_0_90 
* INOUT : bl_0_91 
* INOUT : br_0_91 
* INOUT : bl_0_92 
* INOUT : br_0_92 
* INOUT : bl_0_93 
* INOUT : br_0_93 
* INOUT : bl_0_94 
* INOUT : br_0_94 
* INOUT : bl_0_95 
* INOUT : br_0_95 
* INOUT : bl_0_96 
* INOUT : br_0_96 
* INOUT : bl_0_97 
* INOUT : br_0_97 
* INOUT : bl_0_98 
* INOUT : br_0_98 
* INOUT : bl_0_99 
* INOUT : br_0_99 
* INOUT : bl_0_100 
* INOUT : br_0_100 
* INOUT : bl_0_101 
* INOUT : br_0_101 
* INOUT : bl_0_102 
* INOUT : br_0_102 
* INOUT : bl_0_103 
* INOUT : br_0_103 
* INOUT : bl_0_104 
* INOUT : br_0_104 
* INOUT : bl_0_105 
* INOUT : br_0_105 
* INOUT : bl_0_106 
* INOUT : br_0_106 
* INOUT : bl_0_107 
* INOUT : br_0_107 
* INOUT : bl_0_108 
* INOUT : br_0_108 
* INOUT : bl_0_109 
* INOUT : br_0_109 
* INOUT : bl_0_110 
* INOUT : br_0_110 
* INOUT : bl_0_111 
* INOUT : br_0_111 
* INOUT : bl_0_112 
* INOUT : br_0_112 
* INOUT : bl_0_113 
* INOUT : br_0_113 
* INOUT : bl_0_114 
* INOUT : br_0_114 
* INOUT : bl_0_115 
* INOUT : br_0_115 
* INOUT : bl_0_116 
* INOUT : br_0_116 
* INOUT : bl_0_117 
* INOUT : br_0_117 
* INOUT : bl_0_118 
* INOUT : br_0_118 
* INOUT : bl_0_119 
* INOUT : br_0_119 
* INOUT : bl_0_120 
* INOUT : br_0_120 
* INOUT : bl_0_121 
* INOUT : br_0_121 
* INOUT : bl_0_122 
* INOUT : br_0_122 
* INOUT : bl_0_123 
* INOUT : br_0_123 
* INOUT : bl_0_124 
* INOUT : br_0_124 
* INOUT : bl_0_125 
* INOUT : br_0_125 
* INOUT : bl_0_126 
* INOUT : br_0_126 
* INOUT : bl_0_127 
* INOUT : br_0_127 
* INOUT : bl_0_128 
* INOUT : br_0_128 
* INOUT : bl_0_129 
* INOUT : br_0_129 
* INOUT : bl_0_130 
* INOUT : br_0_130 
* INOUT : bl_0_131 
* INOUT : br_0_131 
* INOUT : bl_0_132 
* INOUT : br_0_132 
* INOUT : bl_0_133 
* INOUT : br_0_133 
* INOUT : bl_0_134 
* INOUT : br_0_134 
* INOUT : bl_0_135 
* INOUT : br_0_135 
* INOUT : bl_0_136 
* INOUT : br_0_136 
* INOUT : bl_0_137 
* INOUT : br_0_137 
* INOUT : bl_0_138 
* INOUT : br_0_138 
* INOUT : bl_0_139 
* INOUT : br_0_139 
* INOUT : bl_0_140 
* INOUT : br_0_140 
* INOUT : bl_0_141 
* INOUT : br_0_141 
* INOUT : bl_0_142 
* INOUT : br_0_142 
* INOUT : bl_0_143 
* INOUT : br_0_143 
* INOUT : bl_0_144 
* INOUT : br_0_144 
* INOUT : bl_0_145 
* INOUT : br_0_145 
* INOUT : bl_0_146 
* INOUT : br_0_146 
* INOUT : bl_0_147 
* INOUT : br_0_147 
* INOUT : bl_0_148 
* INOUT : br_0_148 
* INOUT : bl_0_149 
* INOUT : br_0_149 
* INOUT : bl_0_150 
* INOUT : br_0_150 
* INOUT : bl_0_151 
* INOUT : br_0_151 
* INOUT : bl_0_152 
* INOUT : br_0_152 
* INOUT : bl_0_153 
* INOUT : br_0_153 
* INOUT : bl_0_154 
* INOUT : br_0_154 
* INOUT : bl_0_155 
* INOUT : br_0_155 
* INOUT : bl_0_156 
* INOUT : br_0_156 
* INOUT : bl_0_157 
* INOUT : br_0_157 
* INOUT : bl_0_158 
* INOUT : br_0_158 
* INOUT : bl_0_159 
* INOUT : br_0_159 
* INOUT : bl_0_160 
* INOUT : br_0_160 
* INOUT : bl_0_161 
* INOUT : br_0_161 
* INOUT : bl_0_162 
* INOUT : br_0_162 
* INOUT : bl_0_163 
* INOUT : br_0_163 
* INOUT : bl_0_164 
* INOUT : br_0_164 
* INOUT : bl_0_165 
* INOUT : br_0_165 
* INOUT : bl_0_166 
* INOUT : br_0_166 
* INOUT : bl_0_167 
* INOUT : br_0_167 
* INOUT : bl_0_168 
* INOUT : br_0_168 
* INOUT : bl_0_169 
* INOUT : br_0_169 
* INOUT : bl_0_170 
* INOUT : br_0_170 
* INOUT : bl_0_171 
* INOUT : br_0_171 
* INOUT : bl_0_172 
* INOUT : br_0_172 
* INOUT : bl_0_173 
* INOUT : br_0_173 
* INOUT : bl_0_174 
* INOUT : br_0_174 
* INOUT : bl_0_175 
* INOUT : br_0_175 
* INOUT : bl_0_176 
* INOUT : br_0_176 
* INOUT : bl_0_177 
* INOUT : br_0_177 
* INOUT : bl_0_178 
* INOUT : br_0_178 
* INOUT : bl_0_179 
* INOUT : br_0_179 
* INOUT : bl_0_180 
* INOUT : br_0_180 
* INOUT : bl_0_181 
* INOUT : br_0_181 
* INOUT : bl_0_182 
* INOUT : br_0_182 
* INOUT : bl_0_183 
* INOUT : br_0_183 
* INOUT : bl_0_184 
* INOUT : br_0_184 
* INOUT : bl_0_185 
* INOUT : br_0_185 
* INOUT : bl_0_186 
* INOUT : br_0_186 
* INOUT : bl_0_187 
* INOUT : br_0_187 
* INOUT : bl_0_188 
* INOUT : br_0_188 
* INOUT : bl_0_189 
* INOUT : br_0_189 
* INOUT : bl_0_190 
* INOUT : br_0_190 
* INOUT : bl_0_191 
* INOUT : br_0_191 
* INOUT : bl_0_192 
* INOUT : br_0_192 
* INOUT : bl_0_193 
* INOUT : br_0_193 
* INOUT : bl_0_194 
* INOUT : br_0_194 
* INOUT : bl_0_195 
* INOUT : br_0_195 
* INOUT : bl_0_196 
* INOUT : br_0_196 
* INOUT : bl_0_197 
* INOUT : br_0_197 
* INOUT : bl_0_198 
* INOUT : br_0_198 
* INOUT : bl_0_199 
* INOUT : br_0_199 
* INOUT : bl_0_200 
* INOUT : br_0_200 
* INOUT : bl_0_201 
* INOUT : br_0_201 
* INOUT : bl_0_202 
* INOUT : br_0_202 
* INOUT : bl_0_203 
* INOUT : br_0_203 
* INOUT : bl_0_204 
* INOUT : br_0_204 
* INOUT : bl_0_205 
* INOUT : br_0_205 
* INOUT : bl_0_206 
* INOUT : br_0_206 
* INOUT : bl_0_207 
* INOUT : br_0_207 
* INOUT : bl_0_208 
* INOUT : br_0_208 
* INOUT : bl_0_209 
* INOUT : br_0_209 
* INOUT : bl_0_210 
* INOUT : br_0_210 
* INOUT : bl_0_211 
* INOUT : br_0_211 
* INOUT : bl_0_212 
* INOUT : br_0_212 
* INOUT : bl_0_213 
* INOUT : br_0_213 
* INOUT : bl_0_214 
* INOUT : br_0_214 
* INOUT : bl_0_215 
* INOUT : br_0_215 
* INOUT : bl_0_216 
* INOUT : br_0_216 
* INOUT : bl_0_217 
* INOUT : br_0_217 
* INOUT : bl_0_218 
* INOUT : br_0_218 
* INOUT : bl_0_219 
* INOUT : br_0_219 
* INOUT : bl_0_220 
* INOUT : br_0_220 
* INOUT : bl_0_221 
* INOUT : br_0_221 
* INOUT : bl_0_222 
* INOUT : br_0_222 
* INOUT : bl_0_223 
* INOUT : br_0_223 
* INOUT : bl_0_224 
* INOUT : br_0_224 
* INOUT : bl_0_225 
* INOUT : br_0_225 
* INOUT : bl_0_226 
* INOUT : br_0_226 
* INOUT : bl_0_227 
* INOUT : br_0_227 
* INOUT : bl_0_228 
* INOUT : br_0_228 
* INOUT : bl_0_229 
* INOUT : br_0_229 
* INOUT : bl_0_230 
* INOUT : br_0_230 
* INOUT : bl_0_231 
* INOUT : br_0_231 
* INOUT : bl_0_232 
* INOUT : br_0_232 
* INOUT : bl_0_233 
* INOUT : br_0_233 
* INOUT : bl_0_234 
* INOUT : br_0_234 
* INOUT : bl_0_235 
* INOUT : br_0_235 
* INOUT : bl_0_236 
* INOUT : br_0_236 
* INOUT : bl_0_237 
* INOUT : br_0_237 
* INOUT : bl_0_238 
* INOUT : br_0_238 
* INOUT : bl_0_239 
* INOUT : br_0_239 
* INOUT : bl_0_240 
* INOUT : br_0_240 
* INOUT : bl_0_241 
* INOUT : br_0_241 
* INOUT : bl_0_242 
* INOUT : br_0_242 
* INOUT : bl_0_243 
* INOUT : br_0_243 
* INOUT : bl_0_244 
* INOUT : br_0_244 
* INOUT : bl_0_245 
* INOUT : br_0_245 
* INOUT : bl_0_246 
* INOUT : br_0_246 
* INOUT : bl_0_247 
* INOUT : br_0_247 
* INOUT : bl_0_248 
* INOUT : br_0_248 
* INOUT : bl_0_249 
* INOUT : br_0_249 
* INOUT : bl_0_250 
* INOUT : br_0_250 
* INOUT : bl_0_251 
* INOUT : br_0_251 
* INOUT : bl_0_252 
* INOUT : br_0_252 
* INOUT : bl_0_253 
* INOUT : br_0_253 
* INOUT : bl_0_254 
* INOUT : br_0_254 
* INOUT : bl_0_255 
* INOUT : br_0_255 
* INOUT : bl_0_256 
* INOUT : br_0_256 
* INPUT : wl_0_0 
* POWER : vdd 
* GROUND: gnd 
Xbit_r0_c0
+ bl_0_0 br_0_0 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c1
+ bl_0_1 br_0_1 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c2
+ bl_0_2 br_0_2 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c3
+ bl_0_3 br_0_3 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c4
+ bl_0_4 br_0_4 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c5
+ bl_0_5 br_0_5 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c6
+ bl_0_6 br_0_6 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c7
+ bl_0_7 br_0_7 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c8
+ bl_0_8 br_0_8 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c9
+ bl_0_9 br_0_9 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c10
+ bl_0_10 br_0_10 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c11
+ bl_0_11 br_0_11 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c12
+ bl_0_12 br_0_12 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c13
+ bl_0_13 br_0_13 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c14
+ bl_0_14 br_0_14 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c15
+ bl_0_15 br_0_15 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c16
+ bl_0_16 br_0_16 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c17
+ bl_0_17 br_0_17 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c18
+ bl_0_18 br_0_18 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c19
+ bl_0_19 br_0_19 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c20
+ bl_0_20 br_0_20 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c21
+ bl_0_21 br_0_21 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c22
+ bl_0_22 br_0_22 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c23
+ bl_0_23 br_0_23 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c24
+ bl_0_24 br_0_24 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c25
+ bl_0_25 br_0_25 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c26
+ bl_0_26 br_0_26 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c27
+ bl_0_27 br_0_27 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c28
+ bl_0_28 br_0_28 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c29
+ bl_0_29 br_0_29 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c30
+ bl_0_30 br_0_30 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c31
+ bl_0_31 br_0_31 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c32
+ bl_0_32 br_0_32 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c33
+ bl_0_33 br_0_33 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c34
+ bl_0_34 br_0_34 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c35
+ bl_0_35 br_0_35 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c36
+ bl_0_36 br_0_36 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c37
+ bl_0_37 br_0_37 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c38
+ bl_0_38 br_0_38 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c39
+ bl_0_39 br_0_39 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c40
+ bl_0_40 br_0_40 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c41
+ bl_0_41 br_0_41 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c42
+ bl_0_42 br_0_42 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c43
+ bl_0_43 br_0_43 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c44
+ bl_0_44 br_0_44 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c45
+ bl_0_45 br_0_45 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c46
+ bl_0_46 br_0_46 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c47
+ bl_0_47 br_0_47 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c48
+ bl_0_48 br_0_48 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c49
+ bl_0_49 br_0_49 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c50
+ bl_0_50 br_0_50 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c51
+ bl_0_51 br_0_51 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c52
+ bl_0_52 br_0_52 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c53
+ bl_0_53 br_0_53 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c54
+ bl_0_54 br_0_54 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c55
+ bl_0_55 br_0_55 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c56
+ bl_0_56 br_0_56 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c57
+ bl_0_57 br_0_57 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c58
+ bl_0_58 br_0_58 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c59
+ bl_0_59 br_0_59 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c60
+ bl_0_60 br_0_60 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c61
+ bl_0_61 br_0_61 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c62
+ bl_0_62 br_0_62 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c63
+ bl_0_63 br_0_63 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c64
+ bl_0_64 br_0_64 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c65
+ bl_0_65 br_0_65 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c66
+ bl_0_66 br_0_66 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c67
+ bl_0_67 br_0_67 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c68
+ bl_0_68 br_0_68 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c69
+ bl_0_69 br_0_69 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c70
+ bl_0_70 br_0_70 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c71
+ bl_0_71 br_0_71 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c72
+ bl_0_72 br_0_72 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c73
+ bl_0_73 br_0_73 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c74
+ bl_0_74 br_0_74 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c75
+ bl_0_75 br_0_75 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c76
+ bl_0_76 br_0_76 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c77
+ bl_0_77 br_0_77 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c78
+ bl_0_78 br_0_78 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c79
+ bl_0_79 br_0_79 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c80
+ bl_0_80 br_0_80 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c81
+ bl_0_81 br_0_81 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c82
+ bl_0_82 br_0_82 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c83
+ bl_0_83 br_0_83 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c84
+ bl_0_84 br_0_84 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c85
+ bl_0_85 br_0_85 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c86
+ bl_0_86 br_0_86 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c87
+ bl_0_87 br_0_87 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c88
+ bl_0_88 br_0_88 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c89
+ bl_0_89 br_0_89 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c90
+ bl_0_90 br_0_90 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c91
+ bl_0_91 br_0_91 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c92
+ bl_0_92 br_0_92 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c93
+ bl_0_93 br_0_93 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c94
+ bl_0_94 br_0_94 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c95
+ bl_0_95 br_0_95 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c96
+ bl_0_96 br_0_96 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c97
+ bl_0_97 br_0_97 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c98
+ bl_0_98 br_0_98 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c99
+ bl_0_99 br_0_99 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c100
+ bl_0_100 br_0_100 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c101
+ bl_0_101 br_0_101 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c102
+ bl_0_102 br_0_102 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c103
+ bl_0_103 br_0_103 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c104
+ bl_0_104 br_0_104 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c105
+ bl_0_105 br_0_105 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c106
+ bl_0_106 br_0_106 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c107
+ bl_0_107 br_0_107 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c108
+ bl_0_108 br_0_108 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c109
+ bl_0_109 br_0_109 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c110
+ bl_0_110 br_0_110 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c111
+ bl_0_111 br_0_111 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c112
+ bl_0_112 br_0_112 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c113
+ bl_0_113 br_0_113 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c114
+ bl_0_114 br_0_114 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c115
+ bl_0_115 br_0_115 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c116
+ bl_0_116 br_0_116 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c117
+ bl_0_117 br_0_117 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c118
+ bl_0_118 br_0_118 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c119
+ bl_0_119 br_0_119 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c120
+ bl_0_120 br_0_120 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c121
+ bl_0_121 br_0_121 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c122
+ bl_0_122 br_0_122 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c123
+ bl_0_123 br_0_123 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c124
+ bl_0_124 br_0_124 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c125
+ bl_0_125 br_0_125 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c126
+ bl_0_126 br_0_126 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c127
+ bl_0_127 br_0_127 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c128
+ bl_0_128 br_0_128 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c129
+ bl_0_129 br_0_129 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c130
+ bl_0_130 br_0_130 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c131
+ bl_0_131 br_0_131 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c132
+ bl_0_132 br_0_132 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c133
+ bl_0_133 br_0_133 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c134
+ bl_0_134 br_0_134 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c135
+ bl_0_135 br_0_135 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c136
+ bl_0_136 br_0_136 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c137
+ bl_0_137 br_0_137 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c138
+ bl_0_138 br_0_138 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c139
+ bl_0_139 br_0_139 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c140
+ bl_0_140 br_0_140 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c141
+ bl_0_141 br_0_141 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c142
+ bl_0_142 br_0_142 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c143
+ bl_0_143 br_0_143 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c144
+ bl_0_144 br_0_144 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c145
+ bl_0_145 br_0_145 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c146
+ bl_0_146 br_0_146 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c147
+ bl_0_147 br_0_147 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c148
+ bl_0_148 br_0_148 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c149
+ bl_0_149 br_0_149 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c150
+ bl_0_150 br_0_150 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c151
+ bl_0_151 br_0_151 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c152
+ bl_0_152 br_0_152 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c153
+ bl_0_153 br_0_153 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c154
+ bl_0_154 br_0_154 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c155
+ bl_0_155 br_0_155 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c156
+ bl_0_156 br_0_156 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c157
+ bl_0_157 br_0_157 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c158
+ bl_0_158 br_0_158 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c159
+ bl_0_159 br_0_159 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c160
+ bl_0_160 br_0_160 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c161
+ bl_0_161 br_0_161 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c162
+ bl_0_162 br_0_162 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c163
+ bl_0_163 br_0_163 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c164
+ bl_0_164 br_0_164 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c165
+ bl_0_165 br_0_165 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c166
+ bl_0_166 br_0_166 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c167
+ bl_0_167 br_0_167 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c168
+ bl_0_168 br_0_168 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c169
+ bl_0_169 br_0_169 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c170
+ bl_0_170 br_0_170 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c171
+ bl_0_171 br_0_171 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c172
+ bl_0_172 br_0_172 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c173
+ bl_0_173 br_0_173 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c174
+ bl_0_174 br_0_174 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c175
+ bl_0_175 br_0_175 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c176
+ bl_0_176 br_0_176 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c177
+ bl_0_177 br_0_177 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c178
+ bl_0_178 br_0_178 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c179
+ bl_0_179 br_0_179 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c180
+ bl_0_180 br_0_180 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c181
+ bl_0_181 br_0_181 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c182
+ bl_0_182 br_0_182 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c183
+ bl_0_183 br_0_183 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c184
+ bl_0_184 br_0_184 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c185
+ bl_0_185 br_0_185 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c186
+ bl_0_186 br_0_186 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c187
+ bl_0_187 br_0_187 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c188
+ bl_0_188 br_0_188 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c189
+ bl_0_189 br_0_189 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c190
+ bl_0_190 br_0_190 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c191
+ bl_0_191 br_0_191 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c192
+ bl_0_192 br_0_192 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c193
+ bl_0_193 br_0_193 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c194
+ bl_0_194 br_0_194 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c195
+ bl_0_195 br_0_195 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c196
+ bl_0_196 br_0_196 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c197
+ bl_0_197 br_0_197 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c198
+ bl_0_198 br_0_198 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c199
+ bl_0_199 br_0_199 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c200
+ bl_0_200 br_0_200 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c201
+ bl_0_201 br_0_201 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c202
+ bl_0_202 br_0_202 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c203
+ bl_0_203 br_0_203 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c204
+ bl_0_204 br_0_204 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c205
+ bl_0_205 br_0_205 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c206
+ bl_0_206 br_0_206 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c207
+ bl_0_207 br_0_207 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c208
+ bl_0_208 br_0_208 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c209
+ bl_0_209 br_0_209 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c210
+ bl_0_210 br_0_210 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c211
+ bl_0_211 br_0_211 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c212
+ bl_0_212 br_0_212 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c213
+ bl_0_213 br_0_213 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c214
+ bl_0_214 br_0_214 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c215
+ bl_0_215 br_0_215 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c216
+ bl_0_216 br_0_216 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c217
+ bl_0_217 br_0_217 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c218
+ bl_0_218 br_0_218 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c219
+ bl_0_219 br_0_219 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c220
+ bl_0_220 br_0_220 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c221
+ bl_0_221 br_0_221 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c222
+ bl_0_222 br_0_222 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c223
+ bl_0_223 br_0_223 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c224
+ bl_0_224 br_0_224 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c225
+ bl_0_225 br_0_225 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c226
+ bl_0_226 br_0_226 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c227
+ bl_0_227 br_0_227 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c228
+ bl_0_228 br_0_228 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c229
+ bl_0_229 br_0_229 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c230
+ bl_0_230 br_0_230 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c231
+ bl_0_231 br_0_231 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c232
+ bl_0_232 br_0_232 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c233
+ bl_0_233 br_0_233 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c234
+ bl_0_234 br_0_234 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c235
+ bl_0_235 br_0_235 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c236
+ bl_0_236 br_0_236 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c237
+ bl_0_237 br_0_237 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c238
+ bl_0_238 br_0_238 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c239
+ bl_0_239 br_0_239 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c240
+ bl_0_240 br_0_240 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c241
+ bl_0_241 br_0_241 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c242
+ bl_0_242 br_0_242 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c243
+ bl_0_243 br_0_243 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c244
+ bl_0_244 br_0_244 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c245
+ bl_0_245 br_0_245 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c246
+ bl_0_246 br_0_246 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c247
+ bl_0_247 br_0_247 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c248
+ bl_0_248 br_0_248 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c249
+ bl_0_249 br_0_249 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c250
+ bl_0_250 br_0_250 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c251
+ bl_0_251 br_0_251 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c252
+ bl_0_252 br_0_252 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c253
+ bl_0_253 br_0_253 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c254
+ bl_0_254 br_0_254 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c255
+ bl_0_255 br_0_255 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c256
+ bl_0_256 br_0_256 wl_0_0 vdd gnd
+ dummy_cell_1rw
.ENDS sram_1rw0r0w_32_1024_freepdk45_dummy_array_1

.SUBCKT replica_cell_1rw bl br wl vdd gnd
* Inverter 1
MM0 vdd Q gnd gnd NMOS_VTG W=205.00n L=50n
MM4 vdd Q vdd vdd PMOS_VTG W=90n L=50n

* Inverer 2
MM1 Q vdd gnd gnd NMOS_VTG W=205.00n L=50n
MM5 Q vdd vdd vdd PMOS_VTG W=90n L=50n

* Access transistors
MM3 bl wl Q gnd NMOS_VTG W=135.00n L=50n
MM2 br wl vdd gnd NMOS_VTG W=135.00n L=50n
.ENDS cell_1rw


.SUBCKT sram_1rw0r0w_32_1024_freepdk45_replica_column
+ bl_0_0 br_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7
+ wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16
+ wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24
+ wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32
+ wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40
+ wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48
+ wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56
+ wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64
+ wl_0_65 wl_0_66 wl_0_67 wl_0_68 wl_0_69 wl_0_70 wl_0_71 wl_0_72
+ wl_0_73 wl_0_74 wl_0_75 wl_0_76 wl_0_77 wl_0_78 wl_0_79 wl_0_80
+ wl_0_81 wl_0_82 wl_0_83 wl_0_84 wl_0_85 wl_0_86 wl_0_87 wl_0_88
+ wl_0_89 wl_0_90 wl_0_91 wl_0_92 wl_0_93 wl_0_94 wl_0_95 wl_0_96
+ wl_0_97 wl_0_98 wl_0_99 wl_0_100 wl_0_101 wl_0_102 wl_0_103 wl_0_104
+ wl_0_105 wl_0_106 wl_0_107 wl_0_108 wl_0_109 wl_0_110 wl_0_111
+ wl_0_112 wl_0_113 wl_0_114 wl_0_115 wl_0_116 wl_0_117 wl_0_118
+ wl_0_119 wl_0_120 wl_0_121 wl_0_122 wl_0_123 wl_0_124 wl_0_125
+ wl_0_126 wl_0_127 wl_0_128 vdd gnd
* OUTPUT: bl_0_0 
* OUTPUT: br_0_0 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* INPUT : wl_0_33 
* INPUT : wl_0_34 
* INPUT : wl_0_35 
* INPUT : wl_0_36 
* INPUT : wl_0_37 
* INPUT : wl_0_38 
* INPUT : wl_0_39 
* INPUT : wl_0_40 
* INPUT : wl_0_41 
* INPUT : wl_0_42 
* INPUT : wl_0_43 
* INPUT : wl_0_44 
* INPUT : wl_0_45 
* INPUT : wl_0_46 
* INPUT : wl_0_47 
* INPUT : wl_0_48 
* INPUT : wl_0_49 
* INPUT : wl_0_50 
* INPUT : wl_0_51 
* INPUT : wl_0_52 
* INPUT : wl_0_53 
* INPUT : wl_0_54 
* INPUT : wl_0_55 
* INPUT : wl_0_56 
* INPUT : wl_0_57 
* INPUT : wl_0_58 
* INPUT : wl_0_59 
* INPUT : wl_0_60 
* INPUT : wl_0_61 
* INPUT : wl_0_62 
* INPUT : wl_0_63 
* INPUT : wl_0_64 
* INPUT : wl_0_65 
* INPUT : wl_0_66 
* INPUT : wl_0_67 
* INPUT : wl_0_68 
* INPUT : wl_0_69 
* INPUT : wl_0_70 
* INPUT : wl_0_71 
* INPUT : wl_0_72 
* INPUT : wl_0_73 
* INPUT : wl_0_74 
* INPUT : wl_0_75 
* INPUT : wl_0_76 
* INPUT : wl_0_77 
* INPUT : wl_0_78 
* INPUT : wl_0_79 
* INPUT : wl_0_80 
* INPUT : wl_0_81 
* INPUT : wl_0_82 
* INPUT : wl_0_83 
* INPUT : wl_0_84 
* INPUT : wl_0_85 
* INPUT : wl_0_86 
* INPUT : wl_0_87 
* INPUT : wl_0_88 
* INPUT : wl_0_89 
* INPUT : wl_0_90 
* INPUT : wl_0_91 
* INPUT : wl_0_92 
* INPUT : wl_0_93 
* INPUT : wl_0_94 
* INPUT : wl_0_95 
* INPUT : wl_0_96 
* INPUT : wl_0_97 
* INPUT : wl_0_98 
* INPUT : wl_0_99 
* INPUT : wl_0_100 
* INPUT : wl_0_101 
* INPUT : wl_0_102 
* INPUT : wl_0_103 
* INPUT : wl_0_104 
* INPUT : wl_0_105 
* INPUT : wl_0_106 
* INPUT : wl_0_107 
* INPUT : wl_0_108 
* INPUT : wl_0_109 
* INPUT : wl_0_110 
* INPUT : wl_0_111 
* INPUT : wl_0_112 
* INPUT : wl_0_113 
* INPUT : wl_0_114 
* INPUT : wl_0_115 
* INPUT : wl_0_116 
* INPUT : wl_0_117 
* INPUT : wl_0_118 
* INPUT : wl_0_119 
* INPUT : wl_0_120 
* INPUT : wl_0_121 
* INPUT : wl_0_122 
* INPUT : wl_0_123 
* INPUT : wl_0_124 
* INPUT : wl_0_125 
* INPUT : wl_0_126 
* INPUT : wl_0_127 
* INPUT : wl_0_128 
* POWER : vdd 
* GROUND: gnd 
Xrbc_0
+ bl_0_0 br_0_0 wl_0_0 vdd gnd
+ replica_cell_1rw
Xrbc_1
+ bl_0_0 br_0_0 wl_0_1 vdd gnd
+ replica_cell_1rw
Xrbc_2
+ bl_0_0 br_0_0 wl_0_2 vdd gnd
+ replica_cell_1rw
Xrbc_3
+ bl_0_0 br_0_0 wl_0_3 vdd gnd
+ replica_cell_1rw
Xrbc_4
+ bl_0_0 br_0_0 wl_0_4 vdd gnd
+ replica_cell_1rw
Xrbc_5
+ bl_0_0 br_0_0 wl_0_5 vdd gnd
+ replica_cell_1rw
Xrbc_6
+ bl_0_0 br_0_0 wl_0_6 vdd gnd
+ replica_cell_1rw
Xrbc_7
+ bl_0_0 br_0_0 wl_0_7 vdd gnd
+ replica_cell_1rw
Xrbc_8
+ bl_0_0 br_0_0 wl_0_8 vdd gnd
+ replica_cell_1rw
Xrbc_9
+ bl_0_0 br_0_0 wl_0_9 vdd gnd
+ replica_cell_1rw
Xrbc_10
+ bl_0_0 br_0_0 wl_0_10 vdd gnd
+ replica_cell_1rw
Xrbc_11
+ bl_0_0 br_0_0 wl_0_11 vdd gnd
+ replica_cell_1rw
Xrbc_12
+ bl_0_0 br_0_0 wl_0_12 vdd gnd
+ replica_cell_1rw
Xrbc_13
+ bl_0_0 br_0_0 wl_0_13 vdd gnd
+ replica_cell_1rw
Xrbc_14
+ bl_0_0 br_0_0 wl_0_14 vdd gnd
+ replica_cell_1rw
Xrbc_15
+ bl_0_0 br_0_0 wl_0_15 vdd gnd
+ replica_cell_1rw
Xrbc_16
+ bl_0_0 br_0_0 wl_0_16 vdd gnd
+ replica_cell_1rw
Xrbc_17
+ bl_0_0 br_0_0 wl_0_17 vdd gnd
+ replica_cell_1rw
Xrbc_18
+ bl_0_0 br_0_0 wl_0_18 vdd gnd
+ replica_cell_1rw
Xrbc_19
+ bl_0_0 br_0_0 wl_0_19 vdd gnd
+ replica_cell_1rw
Xrbc_20
+ bl_0_0 br_0_0 wl_0_20 vdd gnd
+ replica_cell_1rw
Xrbc_21
+ bl_0_0 br_0_0 wl_0_21 vdd gnd
+ replica_cell_1rw
Xrbc_22
+ bl_0_0 br_0_0 wl_0_22 vdd gnd
+ replica_cell_1rw
Xrbc_23
+ bl_0_0 br_0_0 wl_0_23 vdd gnd
+ replica_cell_1rw
Xrbc_24
+ bl_0_0 br_0_0 wl_0_24 vdd gnd
+ replica_cell_1rw
Xrbc_25
+ bl_0_0 br_0_0 wl_0_25 vdd gnd
+ replica_cell_1rw
Xrbc_26
+ bl_0_0 br_0_0 wl_0_26 vdd gnd
+ replica_cell_1rw
Xrbc_27
+ bl_0_0 br_0_0 wl_0_27 vdd gnd
+ replica_cell_1rw
Xrbc_28
+ bl_0_0 br_0_0 wl_0_28 vdd gnd
+ replica_cell_1rw
Xrbc_29
+ bl_0_0 br_0_0 wl_0_29 vdd gnd
+ replica_cell_1rw
Xrbc_30
+ bl_0_0 br_0_0 wl_0_30 vdd gnd
+ replica_cell_1rw
Xrbc_31
+ bl_0_0 br_0_0 wl_0_31 vdd gnd
+ replica_cell_1rw
Xrbc_32
+ bl_0_0 br_0_0 wl_0_32 vdd gnd
+ replica_cell_1rw
Xrbc_33
+ bl_0_0 br_0_0 wl_0_33 vdd gnd
+ replica_cell_1rw
Xrbc_34
+ bl_0_0 br_0_0 wl_0_34 vdd gnd
+ replica_cell_1rw
Xrbc_35
+ bl_0_0 br_0_0 wl_0_35 vdd gnd
+ replica_cell_1rw
Xrbc_36
+ bl_0_0 br_0_0 wl_0_36 vdd gnd
+ replica_cell_1rw
Xrbc_37
+ bl_0_0 br_0_0 wl_0_37 vdd gnd
+ replica_cell_1rw
Xrbc_38
+ bl_0_0 br_0_0 wl_0_38 vdd gnd
+ replica_cell_1rw
Xrbc_39
+ bl_0_0 br_0_0 wl_0_39 vdd gnd
+ replica_cell_1rw
Xrbc_40
+ bl_0_0 br_0_0 wl_0_40 vdd gnd
+ replica_cell_1rw
Xrbc_41
+ bl_0_0 br_0_0 wl_0_41 vdd gnd
+ replica_cell_1rw
Xrbc_42
+ bl_0_0 br_0_0 wl_0_42 vdd gnd
+ replica_cell_1rw
Xrbc_43
+ bl_0_0 br_0_0 wl_0_43 vdd gnd
+ replica_cell_1rw
Xrbc_44
+ bl_0_0 br_0_0 wl_0_44 vdd gnd
+ replica_cell_1rw
Xrbc_45
+ bl_0_0 br_0_0 wl_0_45 vdd gnd
+ replica_cell_1rw
Xrbc_46
+ bl_0_0 br_0_0 wl_0_46 vdd gnd
+ replica_cell_1rw
Xrbc_47
+ bl_0_0 br_0_0 wl_0_47 vdd gnd
+ replica_cell_1rw
Xrbc_48
+ bl_0_0 br_0_0 wl_0_48 vdd gnd
+ replica_cell_1rw
Xrbc_49
+ bl_0_0 br_0_0 wl_0_49 vdd gnd
+ replica_cell_1rw
Xrbc_50
+ bl_0_0 br_0_0 wl_0_50 vdd gnd
+ replica_cell_1rw
Xrbc_51
+ bl_0_0 br_0_0 wl_0_51 vdd gnd
+ replica_cell_1rw
Xrbc_52
+ bl_0_0 br_0_0 wl_0_52 vdd gnd
+ replica_cell_1rw
Xrbc_53
+ bl_0_0 br_0_0 wl_0_53 vdd gnd
+ replica_cell_1rw
Xrbc_54
+ bl_0_0 br_0_0 wl_0_54 vdd gnd
+ replica_cell_1rw
Xrbc_55
+ bl_0_0 br_0_0 wl_0_55 vdd gnd
+ replica_cell_1rw
Xrbc_56
+ bl_0_0 br_0_0 wl_0_56 vdd gnd
+ replica_cell_1rw
Xrbc_57
+ bl_0_0 br_0_0 wl_0_57 vdd gnd
+ replica_cell_1rw
Xrbc_58
+ bl_0_0 br_0_0 wl_0_58 vdd gnd
+ replica_cell_1rw
Xrbc_59
+ bl_0_0 br_0_0 wl_0_59 vdd gnd
+ replica_cell_1rw
Xrbc_60
+ bl_0_0 br_0_0 wl_0_60 vdd gnd
+ replica_cell_1rw
Xrbc_61
+ bl_0_0 br_0_0 wl_0_61 vdd gnd
+ replica_cell_1rw
Xrbc_62
+ bl_0_0 br_0_0 wl_0_62 vdd gnd
+ replica_cell_1rw
Xrbc_63
+ bl_0_0 br_0_0 wl_0_63 vdd gnd
+ replica_cell_1rw
Xrbc_64
+ bl_0_0 br_0_0 wl_0_64 vdd gnd
+ replica_cell_1rw
Xrbc_65
+ bl_0_0 br_0_0 wl_0_65 vdd gnd
+ replica_cell_1rw
Xrbc_66
+ bl_0_0 br_0_0 wl_0_66 vdd gnd
+ replica_cell_1rw
Xrbc_67
+ bl_0_0 br_0_0 wl_0_67 vdd gnd
+ replica_cell_1rw
Xrbc_68
+ bl_0_0 br_0_0 wl_0_68 vdd gnd
+ replica_cell_1rw
Xrbc_69
+ bl_0_0 br_0_0 wl_0_69 vdd gnd
+ replica_cell_1rw
Xrbc_70
+ bl_0_0 br_0_0 wl_0_70 vdd gnd
+ replica_cell_1rw
Xrbc_71
+ bl_0_0 br_0_0 wl_0_71 vdd gnd
+ replica_cell_1rw
Xrbc_72
+ bl_0_0 br_0_0 wl_0_72 vdd gnd
+ replica_cell_1rw
Xrbc_73
+ bl_0_0 br_0_0 wl_0_73 vdd gnd
+ replica_cell_1rw
Xrbc_74
+ bl_0_0 br_0_0 wl_0_74 vdd gnd
+ replica_cell_1rw
Xrbc_75
+ bl_0_0 br_0_0 wl_0_75 vdd gnd
+ replica_cell_1rw
Xrbc_76
+ bl_0_0 br_0_0 wl_0_76 vdd gnd
+ replica_cell_1rw
Xrbc_77
+ bl_0_0 br_0_0 wl_0_77 vdd gnd
+ replica_cell_1rw
Xrbc_78
+ bl_0_0 br_0_0 wl_0_78 vdd gnd
+ replica_cell_1rw
Xrbc_79
+ bl_0_0 br_0_0 wl_0_79 vdd gnd
+ replica_cell_1rw
Xrbc_80
+ bl_0_0 br_0_0 wl_0_80 vdd gnd
+ replica_cell_1rw
Xrbc_81
+ bl_0_0 br_0_0 wl_0_81 vdd gnd
+ replica_cell_1rw
Xrbc_82
+ bl_0_0 br_0_0 wl_0_82 vdd gnd
+ replica_cell_1rw
Xrbc_83
+ bl_0_0 br_0_0 wl_0_83 vdd gnd
+ replica_cell_1rw
Xrbc_84
+ bl_0_0 br_0_0 wl_0_84 vdd gnd
+ replica_cell_1rw
Xrbc_85
+ bl_0_0 br_0_0 wl_0_85 vdd gnd
+ replica_cell_1rw
Xrbc_86
+ bl_0_0 br_0_0 wl_0_86 vdd gnd
+ replica_cell_1rw
Xrbc_87
+ bl_0_0 br_0_0 wl_0_87 vdd gnd
+ replica_cell_1rw
Xrbc_88
+ bl_0_0 br_0_0 wl_0_88 vdd gnd
+ replica_cell_1rw
Xrbc_89
+ bl_0_0 br_0_0 wl_0_89 vdd gnd
+ replica_cell_1rw
Xrbc_90
+ bl_0_0 br_0_0 wl_0_90 vdd gnd
+ replica_cell_1rw
Xrbc_91
+ bl_0_0 br_0_0 wl_0_91 vdd gnd
+ replica_cell_1rw
Xrbc_92
+ bl_0_0 br_0_0 wl_0_92 vdd gnd
+ replica_cell_1rw
Xrbc_93
+ bl_0_0 br_0_0 wl_0_93 vdd gnd
+ replica_cell_1rw
Xrbc_94
+ bl_0_0 br_0_0 wl_0_94 vdd gnd
+ replica_cell_1rw
Xrbc_95
+ bl_0_0 br_0_0 wl_0_95 vdd gnd
+ replica_cell_1rw
Xrbc_96
+ bl_0_0 br_0_0 wl_0_96 vdd gnd
+ replica_cell_1rw
Xrbc_97
+ bl_0_0 br_0_0 wl_0_97 vdd gnd
+ replica_cell_1rw
Xrbc_98
+ bl_0_0 br_0_0 wl_0_98 vdd gnd
+ replica_cell_1rw
Xrbc_99
+ bl_0_0 br_0_0 wl_0_99 vdd gnd
+ replica_cell_1rw
Xrbc_100
+ bl_0_0 br_0_0 wl_0_100 vdd gnd
+ replica_cell_1rw
Xrbc_101
+ bl_0_0 br_0_0 wl_0_101 vdd gnd
+ replica_cell_1rw
Xrbc_102
+ bl_0_0 br_0_0 wl_0_102 vdd gnd
+ replica_cell_1rw
Xrbc_103
+ bl_0_0 br_0_0 wl_0_103 vdd gnd
+ replica_cell_1rw
Xrbc_104
+ bl_0_0 br_0_0 wl_0_104 vdd gnd
+ replica_cell_1rw
Xrbc_105
+ bl_0_0 br_0_0 wl_0_105 vdd gnd
+ replica_cell_1rw
Xrbc_106
+ bl_0_0 br_0_0 wl_0_106 vdd gnd
+ replica_cell_1rw
Xrbc_107
+ bl_0_0 br_0_0 wl_0_107 vdd gnd
+ replica_cell_1rw
Xrbc_108
+ bl_0_0 br_0_0 wl_0_108 vdd gnd
+ replica_cell_1rw
Xrbc_109
+ bl_0_0 br_0_0 wl_0_109 vdd gnd
+ replica_cell_1rw
Xrbc_110
+ bl_0_0 br_0_0 wl_0_110 vdd gnd
+ replica_cell_1rw
Xrbc_111
+ bl_0_0 br_0_0 wl_0_111 vdd gnd
+ replica_cell_1rw
Xrbc_112
+ bl_0_0 br_0_0 wl_0_112 vdd gnd
+ replica_cell_1rw
Xrbc_113
+ bl_0_0 br_0_0 wl_0_113 vdd gnd
+ replica_cell_1rw
Xrbc_114
+ bl_0_0 br_0_0 wl_0_114 vdd gnd
+ replica_cell_1rw
Xrbc_115
+ bl_0_0 br_0_0 wl_0_115 vdd gnd
+ replica_cell_1rw
Xrbc_116
+ bl_0_0 br_0_0 wl_0_116 vdd gnd
+ replica_cell_1rw
Xrbc_117
+ bl_0_0 br_0_0 wl_0_117 vdd gnd
+ replica_cell_1rw
Xrbc_118
+ bl_0_0 br_0_0 wl_0_118 vdd gnd
+ replica_cell_1rw
Xrbc_119
+ bl_0_0 br_0_0 wl_0_119 vdd gnd
+ replica_cell_1rw
Xrbc_120
+ bl_0_0 br_0_0 wl_0_120 vdd gnd
+ replica_cell_1rw
Xrbc_121
+ bl_0_0 br_0_0 wl_0_121 vdd gnd
+ replica_cell_1rw
Xrbc_122
+ bl_0_0 br_0_0 wl_0_122 vdd gnd
+ replica_cell_1rw
Xrbc_123
+ bl_0_0 br_0_0 wl_0_123 vdd gnd
+ replica_cell_1rw
Xrbc_124
+ bl_0_0 br_0_0 wl_0_124 vdd gnd
+ replica_cell_1rw
Xrbc_125
+ bl_0_0 br_0_0 wl_0_125 vdd gnd
+ replica_cell_1rw
Xrbc_126
+ bl_0_0 br_0_0 wl_0_126 vdd gnd
+ replica_cell_1rw
Xrbc_127
+ bl_0_0 br_0_0 wl_0_127 vdd gnd
+ replica_cell_1rw
Xrbc_128
+ bl_0_0 br_0_0 wl_0_128 vdd gnd
+ replica_cell_1rw
.ENDS sram_1rw0r0w_32_1024_freepdk45_replica_column

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_dummy_array
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65
+ bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69
+ bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73
+ bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77
+ bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81
+ bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85
+ bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89
+ bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93
+ bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97
+ bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101
+ bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105
+ br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108
+ bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112
+ br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115
+ bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119
+ br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122
+ bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126
+ br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 bl_0_129 br_0_129
+ bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132 br_0_132 bl_0_133
+ br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135 bl_0_136 br_0_136
+ bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139 br_0_139 bl_0_140
+ br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142 bl_0_143 br_0_143
+ bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146 br_0_146 bl_0_147
+ br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149 bl_0_150 br_0_150
+ bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153 br_0_153 bl_0_154
+ br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156 bl_0_157 br_0_157
+ bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160 br_0_160 bl_0_161
+ br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163 bl_0_164 br_0_164
+ bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167 br_0_167 bl_0_168
+ br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170 bl_0_171 br_0_171
+ bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174 br_0_174 bl_0_175
+ br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177 bl_0_178 br_0_178
+ bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181 br_0_181 bl_0_182
+ br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184 bl_0_185 br_0_185
+ bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188 br_0_188 bl_0_189
+ br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191 bl_0_192 br_0_192
+ bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195 br_0_195 bl_0_196
+ br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198 bl_0_199 br_0_199
+ bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202 br_0_202 bl_0_203
+ br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205 bl_0_206 br_0_206
+ bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209 br_0_209 bl_0_210
+ br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212 bl_0_213 br_0_213
+ bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216 br_0_216 bl_0_217
+ br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219 bl_0_220 br_0_220
+ bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223 br_0_223 bl_0_224
+ br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226 bl_0_227 br_0_227
+ bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230 br_0_230 bl_0_231
+ br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233 bl_0_234 br_0_234
+ bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237 br_0_237 bl_0_238
+ br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240 bl_0_241 br_0_241
+ bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244 br_0_244 bl_0_245
+ br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247 bl_0_248 br_0_248
+ bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251 br_0_251 bl_0_252
+ br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254 bl_0_255 br_0_255 wl_0_0
+ vdd gnd
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INOUT : bl_0_64 
* INOUT : br_0_64 
* INOUT : bl_0_65 
* INOUT : br_0_65 
* INOUT : bl_0_66 
* INOUT : br_0_66 
* INOUT : bl_0_67 
* INOUT : br_0_67 
* INOUT : bl_0_68 
* INOUT : br_0_68 
* INOUT : bl_0_69 
* INOUT : br_0_69 
* INOUT : bl_0_70 
* INOUT : br_0_70 
* INOUT : bl_0_71 
* INOUT : br_0_71 
* INOUT : bl_0_72 
* INOUT : br_0_72 
* INOUT : bl_0_73 
* INOUT : br_0_73 
* INOUT : bl_0_74 
* INOUT : br_0_74 
* INOUT : bl_0_75 
* INOUT : br_0_75 
* INOUT : bl_0_76 
* INOUT : br_0_76 
* INOUT : bl_0_77 
* INOUT : br_0_77 
* INOUT : bl_0_78 
* INOUT : br_0_78 
* INOUT : bl_0_79 
* INOUT : br_0_79 
* INOUT : bl_0_80 
* INOUT : br_0_80 
* INOUT : bl_0_81 
* INOUT : br_0_81 
* INOUT : bl_0_82 
* INOUT : br_0_82 
* INOUT : bl_0_83 
* INOUT : br_0_83 
* INOUT : bl_0_84 
* INOUT : br_0_84 
* INOUT : bl_0_85 
* INOUT : br_0_85 
* INOUT : bl_0_86 
* INOUT : br_0_86 
* INOUT : bl_0_87 
* INOUT : br_0_87 
* INOUT : bl_0_88 
* INOUT : br_0_88 
* INOUT : bl_0_89 
* INOUT : br_0_89 
* INOUT : bl_0_90 
* INOUT : br_0_90 
* INOUT : bl_0_91 
* INOUT : br_0_91 
* INOUT : bl_0_92 
* INOUT : br_0_92 
* INOUT : bl_0_93 
* INOUT : br_0_93 
* INOUT : bl_0_94 
* INOUT : br_0_94 
* INOUT : bl_0_95 
* INOUT : br_0_95 
* INOUT : bl_0_96 
* INOUT : br_0_96 
* INOUT : bl_0_97 
* INOUT : br_0_97 
* INOUT : bl_0_98 
* INOUT : br_0_98 
* INOUT : bl_0_99 
* INOUT : br_0_99 
* INOUT : bl_0_100 
* INOUT : br_0_100 
* INOUT : bl_0_101 
* INOUT : br_0_101 
* INOUT : bl_0_102 
* INOUT : br_0_102 
* INOUT : bl_0_103 
* INOUT : br_0_103 
* INOUT : bl_0_104 
* INOUT : br_0_104 
* INOUT : bl_0_105 
* INOUT : br_0_105 
* INOUT : bl_0_106 
* INOUT : br_0_106 
* INOUT : bl_0_107 
* INOUT : br_0_107 
* INOUT : bl_0_108 
* INOUT : br_0_108 
* INOUT : bl_0_109 
* INOUT : br_0_109 
* INOUT : bl_0_110 
* INOUT : br_0_110 
* INOUT : bl_0_111 
* INOUT : br_0_111 
* INOUT : bl_0_112 
* INOUT : br_0_112 
* INOUT : bl_0_113 
* INOUT : br_0_113 
* INOUT : bl_0_114 
* INOUT : br_0_114 
* INOUT : bl_0_115 
* INOUT : br_0_115 
* INOUT : bl_0_116 
* INOUT : br_0_116 
* INOUT : bl_0_117 
* INOUT : br_0_117 
* INOUT : bl_0_118 
* INOUT : br_0_118 
* INOUT : bl_0_119 
* INOUT : br_0_119 
* INOUT : bl_0_120 
* INOUT : br_0_120 
* INOUT : bl_0_121 
* INOUT : br_0_121 
* INOUT : bl_0_122 
* INOUT : br_0_122 
* INOUT : bl_0_123 
* INOUT : br_0_123 
* INOUT : bl_0_124 
* INOUT : br_0_124 
* INOUT : bl_0_125 
* INOUT : br_0_125 
* INOUT : bl_0_126 
* INOUT : br_0_126 
* INOUT : bl_0_127 
* INOUT : br_0_127 
* INOUT : bl_0_128 
* INOUT : br_0_128 
* INOUT : bl_0_129 
* INOUT : br_0_129 
* INOUT : bl_0_130 
* INOUT : br_0_130 
* INOUT : bl_0_131 
* INOUT : br_0_131 
* INOUT : bl_0_132 
* INOUT : br_0_132 
* INOUT : bl_0_133 
* INOUT : br_0_133 
* INOUT : bl_0_134 
* INOUT : br_0_134 
* INOUT : bl_0_135 
* INOUT : br_0_135 
* INOUT : bl_0_136 
* INOUT : br_0_136 
* INOUT : bl_0_137 
* INOUT : br_0_137 
* INOUT : bl_0_138 
* INOUT : br_0_138 
* INOUT : bl_0_139 
* INOUT : br_0_139 
* INOUT : bl_0_140 
* INOUT : br_0_140 
* INOUT : bl_0_141 
* INOUT : br_0_141 
* INOUT : bl_0_142 
* INOUT : br_0_142 
* INOUT : bl_0_143 
* INOUT : br_0_143 
* INOUT : bl_0_144 
* INOUT : br_0_144 
* INOUT : bl_0_145 
* INOUT : br_0_145 
* INOUT : bl_0_146 
* INOUT : br_0_146 
* INOUT : bl_0_147 
* INOUT : br_0_147 
* INOUT : bl_0_148 
* INOUT : br_0_148 
* INOUT : bl_0_149 
* INOUT : br_0_149 
* INOUT : bl_0_150 
* INOUT : br_0_150 
* INOUT : bl_0_151 
* INOUT : br_0_151 
* INOUT : bl_0_152 
* INOUT : br_0_152 
* INOUT : bl_0_153 
* INOUT : br_0_153 
* INOUT : bl_0_154 
* INOUT : br_0_154 
* INOUT : bl_0_155 
* INOUT : br_0_155 
* INOUT : bl_0_156 
* INOUT : br_0_156 
* INOUT : bl_0_157 
* INOUT : br_0_157 
* INOUT : bl_0_158 
* INOUT : br_0_158 
* INOUT : bl_0_159 
* INOUT : br_0_159 
* INOUT : bl_0_160 
* INOUT : br_0_160 
* INOUT : bl_0_161 
* INOUT : br_0_161 
* INOUT : bl_0_162 
* INOUT : br_0_162 
* INOUT : bl_0_163 
* INOUT : br_0_163 
* INOUT : bl_0_164 
* INOUT : br_0_164 
* INOUT : bl_0_165 
* INOUT : br_0_165 
* INOUT : bl_0_166 
* INOUT : br_0_166 
* INOUT : bl_0_167 
* INOUT : br_0_167 
* INOUT : bl_0_168 
* INOUT : br_0_168 
* INOUT : bl_0_169 
* INOUT : br_0_169 
* INOUT : bl_0_170 
* INOUT : br_0_170 
* INOUT : bl_0_171 
* INOUT : br_0_171 
* INOUT : bl_0_172 
* INOUT : br_0_172 
* INOUT : bl_0_173 
* INOUT : br_0_173 
* INOUT : bl_0_174 
* INOUT : br_0_174 
* INOUT : bl_0_175 
* INOUT : br_0_175 
* INOUT : bl_0_176 
* INOUT : br_0_176 
* INOUT : bl_0_177 
* INOUT : br_0_177 
* INOUT : bl_0_178 
* INOUT : br_0_178 
* INOUT : bl_0_179 
* INOUT : br_0_179 
* INOUT : bl_0_180 
* INOUT : br_0_180 
* INOUT : bl_0_181 
* INOUT : br_0_181 
* INOUT : bl_0_182 
* INOUT : br_0_182 
* INOUT : bl_0_183 
* INOUT : br_0_183 
* INOUT : bl_0_184 
* INOUT : br_0_184 
* INOUT : bl_0_185 
* INOUT : br_0_185 
* INOUT : bl_0_186 
* INOUT : br_0_186 
* INOUT : bl_0_187 
* INOUT : br_0_187 
* INOUT : bl_0_188 
* INOUT : br_0_188 
* INOUT : bl_0_189 
* INOUT : br_0_189 
* INOUT : bl_0_190 
* INOUT : br_0_190 
* INOUT : bl_0_191 
* INOUT : br_0_191 
* INOUT : bl_0_192 
* INOUT : br_0_192 
* INOUT : bl_0_193 
* INOUT : br_0_193 
* INOUT : bl_0_194 
* INOUT : br_0_194 
* INOUT : bl_0_195 
* INOUT : br_0_195 
* INOUT : bl_0_196 
* INOUT : br_0_196 
* INOUT : bl_0_197 
* INOUT : br_0_197 
* INOUT : bl_0_198 
* INOUT : br_0_198 
* INOUT : bl_0_199 
* INOUT : br_0_199 
* INOUT : bl_0_200 
* INOUT : br_0_200 
* INOUT : bl_0_201 
* INOUT : br_0_201 
* INOUT : bl_0_202 
* INOUT : br_0_202 
* INOUT : bl_0_203 
* INOUT : br_0_203 
* INOUT : bl_0_204 
* INOUT : br_0_204 
* INOUT : bl_0_205 
* INOUT : br_0_205 
* INOUT : bl_0_206 
* INOUT : br_0_206 
* INOUT : bl_0_207 
* INOUT : br_0_207 
* INOUT : bl_0_208 
* INOUT : br_0_208 
* INOUT : bl_0_209 
* INOUT : br_0_209 
* INOUT : bl_0_210 
* INOUT : br_0_210 
* INOUT : bl_0_211 
* INOUT : br_0_211 
* INOUT : bl_0_212 
* INOUT : br_0_212 
* INOUT : bl_0_213 
* INOUT : br_0_213 
* INOUT : bl_0_214 
* INOUT : br_0_214 
* INOUT : bl_0_215 
* INOUT : br_0_215 
* INOUT : bl_0_216 
* INOUT : br_0_216 
* INOUT : bl_0_217 
* INOUT : br_0_217 
* INOUT : bl_0_218 
* INOUT : br_0_218 
* INOUT : bl_0_219 
* INOUT : br_0_219 
* INOUT : bl_0_220 
* INOUT : br_0_220 
* INOUT : bl_0_221 
* INOUT : br_0_221 
* INOUT : bl_0_222 
* INOUT : br_0_222 
* INOUT : bl_0_223 
* INOUT : br_0_223 
* INOUT : bl_0_224 
* INOUT : br_0_224 
* INOUT : bl_0_225 
* INOUT : br_0_225 
* INOUT : bl_0_226 
* INOUT : br_0_226 
* INOUT : bl_0_227 
* INOUT : br_0_227 
* INOUT : bl_0_228 
* INOUT : br_0_228 
* INOUT : bl_0_229 
* INOUT : br_0_229 
* INOUT : bl_0_230 
* INOUT : br_0_230 
* INOUT : bl_0_231 
* INOUT : br_0_231 
* INOUT : bl_0_232 
* INOUT : br_0_232 
* INOUT : bl_0_233 
* INOUT : br_0_233 
* INOUT : bl_0_234 
* INOUT : br_0_234 
* INOUT : bl_0_235 
* INOUT : br_0_235 
* INOUT : bl_0_236 
* INOUT : br_0_236 
* INOUT : bl_0_237 
* INOUT : br_0_237 
* INOUT : bl_0_238 
* INOUT : br_0_238 
* INOUT : bl_0_239 
* INOUT : br_0_239 
* INOUT : bl_0_240 
* INOUT : br_0_240 
* INOUT : bl_0_241 
* INOUT : br_0_241 
* INOUT : bl_0_242 
* INOUT : br_0_242 
* INOUT : bl_0_243 
* INOUT : br_0_243 
* INOUT : bl_0_244 
* INOUT : br_0_244 
* INOUT : bl_0_245 
* INOUT : br_0_245 
* INOUT : bl_0_246 
* INOUT : br_0_246 
* INOUT : bl_0_247 
* INOUT : br_0_247 
* INOUT : bl_0_248 
* INOUT : br_0_248 
* INOUT : bl_0_249 
* INOUT : br_0_249 
* INOUT : bl_0_250 
* INOUT : br_0_250 
* INOUT : bl_0_251 
* INOUT : br_0_251 
* INOUT : bl_0_252 
* INOUT : br_0_252 
* INOUT : bl_0_253 
* INOUT : br_0_253 
* INOUT : bl_0_254 
* INOUT : br_0_254 
* INOUT : bl_0_255 
* INOUT : br_0_255 
* INPUT : wl_0_0 
* POWER : vdd 
* GROUND: gnd 
Xbit_r0_c0
+ bl_0_0 br_0_0 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c1
+ bl_0_1 br_0_1 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c2
+ bl_0_2 br_0_2 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c3
+ bl_0_3 br_0_3 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c4
+ bl_0_4 br_0_4 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c5
+ bl_0_5 br_0_5 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c6
+ bl_0_6 br_0_6 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c7
+ bl_0_7 br_0_7 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c8
+ bl_0_8 br_0_8 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c9
+ bl_0_9 br_0_9 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c10
+ bl_0_10 br_0_10 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c11
+ bl_0_11 br_0_11 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c12
+ bl_0_12 br_0_12 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c13
+ bl_0_13 br_0_13 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c14
+ bl_0_14 br_0_14 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c15
+ bl_0_15 br_0_15 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c16
+ bl_0_16 br_0_16 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c17
+ bl_0_17 br_0_17 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c18
+ bl_0_18 br_0_18 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c19
+ bl_0_19 br_0_19 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c20
+ bl_0_20 br_0_20 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c21
+ bl_0_21 br_0_21 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c22
+ bl_0_22 br_0_22 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c23
+ bl_0_23 br_0_23 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c24
+ bl_0_24 br_0_24 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c25
+ bl_0_25 br_0_25 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c26
+ bl_0_26 br_0_26 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c27
+ bl_0_27 br_0_27 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c28
+ bl_0_28 br_0_28 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c29
+ bl_0_29 br_0_29 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c30
+ bl_0_30 br_0_30 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c31
+ bl_0_31 br_0_31 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c32
+ bl_0_32 br_0_32 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c33
+ bl_0_33 br_0_33 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c34
+ bl_0_34 br_0_34 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c35
+ bl_0_35 br_0_35 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c36
+ bl_0_36 br_0_36 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c37
+ bl_0_37 br_0_37 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c38
+ bl_0_38 br_0_38 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c39
+ bl_0_39 br_0_39 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c40
+ bl_0_40 br_0_40 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c41
+ bl_0_41 br_0_41 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c42
+ bl_0_42 br_0_42 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c43
+ bl_0_43 br_0_43 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c44
+ bl_0_44 br_0_44 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c45
+ bl_0_45 br_0_45 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c46
+ bl_0_46 br_0_46 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c47
+ bl_0_47 br_0_47 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c48
+ bl_0_48 br_0_48 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c49
+ bl_0_49 br_0_49 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c50
+ bl_0_50 br_0_50 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c51
+ bl_0_51 br_0_51 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c52
+ bl_0_52 br_0_52 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c53
+ bl_0_53 br_0_53 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c54
+ bl_0_54 br_0_54 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c55
+ bl_0_55 br_0_55 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c56
+ bl_0_56 br_0_56 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c57
+ bl_0_57 br_0_57 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c58
+ bl_0_58 br_0_58 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c59
+ bl_0_59 br_0_59 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c60
+ bl_0_60 br_0_60 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c61
+ bl_0_61 br_0_61 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c62
+ bl_0_62 br_0_62 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c63
+ bl_0_63 br_0_63 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c64
+ bl_0_64 br_0_64 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c65
+ bl_0_65 br_0_65 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c66
+ bl_0_66 br_0_66 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c67
+ bl_0_67 br_0_67 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c68
+ bl_0_68 br_0_68 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c69
+ bl_0_69 br_0_69 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c70
+ bl_0_70 br_0_70 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c71
+ bl_0_71 br_0_71 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c72
+ bl_0_72 br_0_72 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c73
+ bl_0_73 br_0_73 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c74
+ bl_0_74 br_0_74 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c75
+ bl_0_75 br_0_75 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c76
+ bl_0_76 br_0_76 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c77
+ bl_0_77 br_0_77 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c78
+ bl_0_78 br_0_78 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c79
+ bl_0_79 br_0_79 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c80
+ bl_0_80 br_0_80 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c81
+ bl_0_81 br_0_81 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c82
+ bl_0_82 br_0_82 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c83
+ bl_0_83 br_0_83 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c84
+ bl_0_84 br_0_84 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c85
+ bl_0_85 br_0_85 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c86
+ bl_0_86 br_0_86 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c87
+ bl_0_87 br_0_87 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c88
+ bl_0_88 br_0_88 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c89
+ bl_0_89 br_0_89 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c90
+ bl_0_90 br_0_90 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c91
+ bl_0_91 br_0_91 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c92
+ bl_0_92 br_0_92 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c93
+ bl_0_93 br_0_93 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c94
+ bl_0_94 br_0_94 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c95
+ bl_0_95 br_0_95 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c96
+ bl_0_96 br_0_96 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c97
+ bl_0_97 br_0_97 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c98
+ bl_0_98 br_0_98 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c99
+ bl_0_99 br_0_99 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c100
+ bl_0_100 br_0_100 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c101
+ bl_0_101 br_0_101 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c102
+ bl_0_102 br_0_102 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c103
+ bl_0_103 br_0_103 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c104
+ bl_0_104 br_0_104 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c105
+ bl_0_105 br_0_105 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c106
+ bl_0_106 br_0_106 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c107
+ bl_0_107 br_0_107 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c108
+ bl_0_108 br_0_108 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c109
+ bl_0_109 br_0_109 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c110
+ bl_0_110 br_0_110 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c111
+ bl_0_111 br_0_111 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c112
+ bl_0_112 br_0_112 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c113
+ bl_0_113 br_0_113 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c114
+ bl_0_114 br_0_114 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c115
+ bl_0_115 br_0_115 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c116
+ bl_0_116 br_0_116 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c117
+ bl_0_117 br_0_117 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c118
+ bl_0_118 br_0_118 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c119
+ bl_0_119 br_0_119 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c120
+ bl_0_120 br_0_120 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c121
+ bl_0_121 br_0_121 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c122
+ bl_0_122 br_0_122 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c123
+ bl_0_123 br_0_123 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c124
+ bl_0_124 br_0_124 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c125
+ bl_0_125 br_0_125 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c126
+ bl_0_126 br_0_126 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c127
+ bl_0_127 br_0_127 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c128
+ bl_0_128 br_0_128 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c129
+ bl_0_129 br_0_129 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c130
+ bl_0_130 br_0_130 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c131
+ bl_0_131 br_0_131 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c132
+ bl_0_132 br_0_132 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c133
+ bl_0_133 br_0_133 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c134
+ bl_0_134 br_0_134 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c135
+ bl_0_135 br_0_135 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c136
+ bl_0_136 br_0_136 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c137
+ bl_0_137 br_0_137 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c138
+ bl_0_138 br_0_138 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c139
+ bl_0_139 br_0_139 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c140
+ bl_0_140 br_0_140 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c141
+ bl_0_141 br_0_141 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c142
+ bl_0_142 br_0_142 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c143
+ bl_0_143 br_0_143 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c144
+ bl_0_144 br_0_144 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c145
+ bl_0_145 br_0_145 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c146
+ bl_0_146 br_0_146 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c147
+ bl_0_147 br_0_147 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c148
+ bl_0_148 br_0_148 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c149
+ bl_0_149 br_0_149 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c150
+ bl_0_150 br_0_150 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c151
+ bl_0_151 br_0_151 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c152
+ bl_0_152 br_0_152 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c153
+ bl_0_153 br_0_153 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c154
+ bl_0_154 br_0_154 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c155
+ bl_0_155 br_0_155 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c156
+ bl_0_156 br_0_156 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c157
+ bl_0_157 br_0_157 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c158
+ bl_0_158 br_0_158 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c159
+ bl_0_159 br_0_159 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c160
+ bl_0_160 br_0_160 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c161
+ bl_0_161 br_0_161 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c162
+ bl_0_162 br_0_162 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c163
+ bl_0_163 br_0_163 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c164
+ bl_0_164 br_0_164 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c165
+ bl_0_165 br_0_165 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c166
+ bl_0_166 br_0_166 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c167
+ bl_0_167 br_0_167 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c168
+ bl_0_168 br_0_168 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c169
+ bl_0_169 br_0_169 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c170
+ bl_0_170 br_0_170 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c171
+ bl_0_171 br_0_171 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c172
+ bl_0_172 br_0_172 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c173
+ bl_0_173 br_0_173 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c174
+ bl_0_174 br_0_174 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c175
+ bl_0_175 br_0_175 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c176
+ bl_0_176 br_0_176 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c177
+ bl_0_177 br_0_177 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c178
+ bl_0_178 br_0_178 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c179
+ bl_0_179 br_0_179 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c180
+ bl_0_180 br_0_180 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c181
+ bl_0_181 br_0_181 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c182
+ bl_0_182 br_0_182 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c183
+ bl_0_183 br_0_183 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c184
+ bl_0_184 br_0_184 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c185
+ bl_0_185 br_0_185 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c186
+ bl_0_186 br_0_186 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c187
+ bl_0_187 br_0_187 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c188
+ bl_0_188 br_0_188 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c189
+ bl_0_189 br_0_189 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c190
+ bl_0_190 br_0_190 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c191
+ bl_0_191 br_0_191 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c192
+ bl_0_192 br_0_192 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c193
+ bl_0_193 br_0_193 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c194
+ bl_0_194 br_0_194 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c195
+ bl_0_195 br_0_195 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c196
+ bl_0_196 br_0_196 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c197
+ bl_0_197 br_0_197 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c198
+ bl_0_198 br_0_198 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c199
+ bl_0_199 br_0_199 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c200
+ bl_0_200 br_0_200 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c201
+ bl_0_201 br_0_201 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c202
+ bl_0_202 br_0_202 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c203
+ bl_0_203 br_0_203 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c204
+ bl_0_204 br_0_204 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c205
+ bl_0_205 br_0_205 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c206
+ bl_0_206 br_0_206 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c207
+ bl_0_207 br_0_207 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c208
+ bl_0_208 br_0_208 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c209
+ bl_0_209 br_0_209 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c210
+ bl_0_210 br_0_210 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c211
+ bl_0_211 br_0_211 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c212
+ bl_0_212 br_0_212 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c213
+ bl_0_213 br_0_213 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c214
+ bl_0_214 br_0_214 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c215
+ bl_0_215 br_0_215 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c216
+ bl_0_216 br_0_216 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c217
+ bl_0_217 br_0_217 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c218
+ bl_0_218 br_0_218 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c219
+ bl_0_219 br_0_219 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c220
+ bl_0_220 br_0_220 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c221
+ bl_0_221 br_0_221 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c222
+ bl_0_222 br_0_222 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c223
+ bl_0_223 br_0_223 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c224
+ bl_0_224 br_0_224 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c225
+ bl_0_225 br_0_225 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c226
+ bl_0_226 br_0_226 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c227
+ bl_0_227 br_0_227 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c228
+ bl_0_228 br_0_228 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c229
+ bl_0_229 br_0_229 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c230
+ bl_0_230 br_0_230 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c231
+ bl_0_231 br_0_231 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c232
+ bl_0_232 br_0_232 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c233
+ bl_0_233 br_0_233 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c234
+ bl_0_234 br_0_234 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c235
+ bl_0_235 br_0_235 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c236
+ bl_0_236 br_0_236 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c237
+ bl_0_237 br_0_237 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c238
+ bl_0_238 br_0_238 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c239
+ bl_0_239 br_0_239 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c240
+ bl_0_240 br_0_240 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c241
+ bl_0_241 br_0_241 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c242
+ bl_0_242 br_0_242 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c243
+ bl_0_243 br_0_243 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c244
+ bl_0_244 br_0_244 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c245
+ bl_0_245 br_0_245 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c246
+ bl_0_246 br_0_246 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c247
+ bl_0_247 br_0_247 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c248
+ bl_0_248 br_0_248 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c249
+ bl_0_249 br_0_249 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c250
+ bl_0_250 br_0_250 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c251
+ bl_0_251 br_0_251 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c252
+ bl_0_252 br_0_252 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c253
+ bl_0_253 br_0_253 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c254
+ bl_0_254 br_0_254 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c255
+ bl_0_255 br_0_255 wl_0_0 vdd gnd
+ dummy_cell_1rw
.ENDS sram_1rw0r0w_32_1024_freepdk45_dummy_array

.SUBCKT cell_1rw bl br wl vdd gnd
* Inverter 1
MM0 Q_bar Q gnd gnd NMOS_VTG W=205.00n L=50n
MM4 Q_bar Q vdd vdd PMOS_VTG W=90n L=50n

* Inverer 2
MM1 Q Q_bar gnd gnd NMOS_VTG W=205.00n L=50n
MM5 Q Q_bar vdd vdd PMOS_VTG W=90n L=50n

* Access transistors
MM3 bl wl Q gnd NMOS_VTG W=135.00n L=50n
MM2 br wl Q_bar gnd NMOS_VTG W=135.00n L=50n
.ENDS cell_1rw


.SUBCKT sram_1rw0r0w_32_1024_freepdk45_bitcell_array
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65
+ bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69
+ bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73
+ bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77
+ bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81
+ bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85
+ bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89
+ bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93
+ bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97
+ bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101
+ bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105
+ br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108
+ bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112
+ br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115
+ bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119
+ br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122
+ bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126
+ br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 bl_0_129 br_0_129
+ bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132 br_0_132 bl_0_133
+ br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135 bl_0_136 br_0_136
+ bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139 br_0_139 bl_0_140
+ br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142 bl_0_143 br_0_143
+ bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146 br_0_146 bl_0_147
+ br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149 bl_0_150 br_0_150
+ bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153 br_0_153 bl_0_154
+ br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156 bl_0_157 br_0_157
+ bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160 br_0_160 bl_0_161
+ br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163 bl_0_164 br_0_164
+ bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167 br_0_167 bl_0_168
+ br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170 bl_0_171 br_0_171
+ bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174 br_0_174 bl_0_175
+ br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177 bl_0_178 br_0_178
+ bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181 br_0_181 bl_0_182
+ br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184 bl_0_185 br_0_185
+ bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188 br_0_188 bl_0_189
+ br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191 bl_0_192 br_0_192
+ bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195 br_0_195 bl_0_196
+ br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198 bl_0_199 br_0_199
+ bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202 br_0_202 bl_0_203
+ br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205 bl_0_206 br_0_206
+ bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209 br_0_209 bl_0_210
+ br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212 bl_0_213 br_0_213
+ bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216 br_0_216 bl_0_217
+ br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219 bl_0_220 br_0_220
+ bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223 br_0_223 bl_0_224
+ br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226 bl_0_227 br_0_227
+ bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230 br_0_230 bl_0_231
+ br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233 bl_0_234 br_0_234
+ bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237 br_0_237 bl_0_238
+ br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240 bl_0_241 br_0_241
+ bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244 br_0_244 bl_0_245
+ br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247 bl_0_248 br_0_248
+ bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251 br_0_251 bl_0_252
+ br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254 bl_0_255 br_0_255 wl_0_0
+ wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10
+ wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18
+ wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26
+ wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34
+ wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42
+ wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50
+ wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57 wl_0_58
+ wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 wl_0_65 wl_0_66
+ wl_0_67 wl_0_68 wl_0_69 wl_0_70 wl_0_71 wl_0_72 wl_0_73 wl_0_74
+ wl_0_75 wl_0_76 wl_0_77 wl_0_78 wl_0_79 wl_0_80 wl_0_81 wl_0_82
+ wl_0_83 wl_0_84 wl_0_85 wl_0_86 wl_0_87 wl_0_88 wl_0_89 wl_0_90
+ wl_0_91 wl_0_92 wl_0_93 wl_0_94 wl_0_95 wl_0_96 wl_0_97 wl_0_98
+ wl_0_99 wl_0_100 wl_0_101 wl_0_102 wl_0_103 wl_0_104 wl_0_105 wl_0_106
+ wl_0_107 wl_0_108 wl_0_109 wl_0_110 wl_0_111 wl_0_112 wl_0_113
+ wl_0_114 wl_0_115 wl_0_116 wl_0_117 wl_0_118 wl_0_119 wl_0_120
+ wl_0_121 wl_0_122 wl_0_123 wl_0_124 wl_0_125 wl_0_126 wl_0_127 vdd gnd
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INOUT : bl_0_64 
* INOUT : br_0_64 
* INOUT : bl_0_65 
* INOUT : br_0_65 
* INOUT : bl_0_66 
* INOUT : br_0_66 
* INOUT : bl_0_67 
* INOUT : br_0_67 
* INOUT : bl_0_68 
* INOUT : br_0_68 
* INOUT : bl_0_69 
* INOUT : br_0_69 
* INOUT : bl_0_70 
* INOUT : br_0_70 
* INOUT : bl_0_71 
* INOUT : br_0_71 
* INOUT : bl_0_72 
* INOUT : br_0_72 
* INOUT : bl_0_73 
* INOUT : br_0_73 
* INOUT : bl_0_74 
* INOUT : br_0_74 
* INOUT : bl_0_75 
* INOUT : br_0_75 
* INOUT : bl_0_76 
* INOUT : br_0_76 
* INOUT : bl_0_77 
* INOUT : br_0_77 
* INOUT : bl_0_78 
* INOUT : br_0_78 
* INOUT : bl_0_79 
* INOUT : br_0_79 
* INOUT : bl_0_80 
* INOUT : br_0_80 
* INOUT : bl_0_81 
* INOUT : br_0_81 
* INOUT : bl_0_82 
* INOUT : br_0_82 
* INOUT : bl_0_83 
* INOUT : br_0_83 
* INOUT : bl_0_84 
* INOUT : br_0_84 
* INOUT : bl_0_85 
* INOUT : br_0_85 
* INOUT : bl_0_86 
* INOUT : br_0_86 
* INOUT : bl_0_87 
* INOUT : br_0_87 
* INOUT : bl_0_88 
* INOUT : br_0_88 
* INOUT : bl_0_89 
* INOUT : br_0_89 
* INOUT : bl_0_90 
* INOUT : br_0_90 
* INOUT : bl_0_91 
* INOUT : br_0_91 
* INOUT : bl_0_92 
* INOUT : br_0_92 
* INOUT : bl_0_93 
* INOUT : br_0_93 
* INOUT : bl_0_94 
* INOUT : br_0_94 
* INOUT : bl_0_95 
* INOUT : br_0_95 
* INOUT : bl_0_96 
* INOUT : br_0_96 
* INOUT : bl_0_97 
* INOUT : br_0_97 
* INOUT : bl_0_98 
* INOUT : br_0_98 
* INOUT : bl_0_99 
* INOUT : br_0_99 
* INOUT : bl_0_100 
* INOUT : br_0_100 
* INOUT : bl_0_101 
* INOUT : br_0_101 
* INOUT : bl_0_102 
* INOUT : br_0_102 
* INOUT : bl_0_103 
* INOUT : br_0_103 
* INOUT : bl_0_104 
* INOUT : br_0_104 
* INOUT : bl_0_105 
* INOUT : br_0_105 
* INOUT : bl_0_106 
* INOUT : br_0_106 
* INOUT : bl_0_107 
* INOUT : br_0_107 
* INOUT : bl_0_108 
* INOUT : br_0_108 
* INOUT : bl_0_109 
* INOUT : br_0_109 
* INOUT : bl_0_110 
* INOUT : br_0_110 
* INOUT : bl_0_111 
* INOUT : br_0_111 
* INOUT : bl_0_112 
* INOUT : br_0_112 
* INOUT : bl_0_113 
* INOUT : br_0_113 
* INOUT : bl_0_114 
* INOUT : br_0_114 
* INOUT : bl_0_115 
* INOUT : br_0_115 
* INOUT : bl_0_116 
* INOUT : br_0_116 
* INOUT : bl_0_117 
* INOUT : br_0_117 
* INOUT : bl_0_118 
* INOUT : br_0_118 
* INOUT : bl_0_119 
* INOUT : br_0_119 
* INOUT : bl_0_120 
* INOUT : br_0_120 
* INOUT : bl_0_121 
* INOUT : br_0_121 
* INOUT : bl_0_122 
* INOUT : br_0_122 
* INOUT : bl_0_123 
* INOUT : br_0_123 
* INOUT : bl_0_124 
* INOUT : br_0_124 
* INOUT : bl_0_125 
* INOUT : br_0_125 
* INOUT : bl_0_126 
* INOUT : br_0_126 
* INOUT : bl_0_127 
* INOUT : br_0_127 
* INOUT : bl_0_128 
* INOUT : br_0_128 
* INOUT : bl_0_129 
* INOUT : br_0_129 
* INOUT : bl_0_130 
* INOUT : br_0_130 
* INOUT : bl_0_131 
* INOUT : br_0_131 
* INOUT : bl_0_132 
* INOUT : br_0_132 
* INOUT : bl_0_133 
* INOUT : br_0_133 
* INOUT : bl_0_134 
* INOUT : br_0_134 
* INOUT : bl_0_135 
* INOUT : br_0_135 
* INOUT : bl_0_136 
* INOUT : br_0_136 
* INOUT : bl_0_137 
* INOUT : br_0_137 
* INOUT : bl_0_138 
* INOUT : br_0_138 
* INOUT : bl_0_139 
* INOUT : br_0_139 
* INOUT : bl_0_140 
* INOUT : br_0_140 
* INOUT : bl_0_141 
* INOUT : br_0_141 
* INOUT : bl_0_142 
* INOUT : br_0_142 
* INOUT : bl_0_143 
* INOUT : br_0_143 
* INOUT : bl_0_144 
* INOUT : br_0_144 
* INOUT : bl_0_145 
* INOUT : br_0_145 
* INOUT : bl_0_146 
* INOUT : br_0_146 
* INOUT : bl_0_147 
* INOUT : br_0_147 
* INOUT : bl_0_148 
* INOUT : br_0_148 
* INOUT : bl_0_149 
* INOUT : br_0_149 
* INOUT : bl_0_150 
* INOUT : br_0_150 
* INOUT : bl_0_151 
* INOUT : br_0_151 
* INOUT : bl_0_152 
* INOUT : br_0_152 
* INOUT : bl_0_153 
* INOUT : br_0_153 
* INOUT : bl_0_154 
* INOUT : br_0_154 
* INOUT : bl_0_155 
* INOUT : br_0_155 
* INOUT : bl_0_156 
* INOUT : br_0_156 
* INOUT : bl_0_157 
* INOUT : br_0_157 
* INOUT : bl_0_158 
* INOUT : br_0_158 
* INOUT : bl_0_159 
* INOUT : br_0_159 
* INOUT : bl_0_160 
* INOUT : br_0_160 
* INOUT : bl_0_161 
* INOUT : br_0_161 
* INOUT : bl_0_162 
* INOUT : br_0_162 
* INOUT : bl_0_163 
* INOUT : br_0_163 
* INOUT : bl_0_164 
* INOUT : br_0_164 
* INOUT : bl_0_165 
* INOUT : br_0_165 
* INOUT : bl_0_166 
* INOUT : br_0_166 
* INOUT : bl_0_167 
* INOUT : br_0_167 
* INOUT : bl_0_168 
* INOUT : br_0_168 
* INOUT : bl_0_169 
* INOUT : br_0_169 
* INOUT : bl_0_170 
* INOUT : br_0_170 
* INOUT : bl_0_171 
* INOUT : br_0_171 
* INOUT : bl_0_172 
* INOUT : br_0_172 
* INOUT : bl_0_173 
* INOUT : br_0_173 
* INOUT : bl_0_174 
* INOUT : br_0_174 
* INOUT : bl_0_175 
* INOUT : br_0_175 
* INOUT : bl_0_176 
* INOUT : br_0_176 
* INOUT : bl_0_177 
* INOUT : br_0_177 
* INOUT : bl_0_178 
* INOUT : br_0_178 
* INOUT : bl_0_179 
* INOUT : br_0_179 
* INOUT : bl_0_180 
* INOUT : br_0_180 
* INOUT : bl_0_181 
* INOUT : br_0_181 
* INOUT : bl_0_182 
* INOUT : br_0_182 
* INOUT : bl_0_183 
* INOUT : br_0_183 
* INOUT : bl_0_184 
* INOUT : br_0_184 
* INOUT : bl_0_185 
* INOUT : br_0_185 
* INOUT : bl_0_186 
* INOUT : br_0_186 
* INOUT : bl_0_187 
* INOUT : br_0_187 
* INOUT : bl_0_188 
* INOUT : br_0_188 
* INOUT : bl_0_189 
* INOUT : br_0_189 
* INOUT : bl_0_190 
* INOUT : br_0_190 
* INOUT : bl_0_191 
* INOUT : br_0_191 
* INOUT : bl_0_192 
* INOUT : br_0_192 
* INOUT : bl_0_193 
* INOUT : br_0_193 
* INOUT : bl_0_194 
* INOUT : br_0_194 
* INOUT : bl_0_195 
* INOUT : br_0_195 
* INOUT : bl_0_196 
* INOUT : br_0_196 
* INOUT : bl_0_197 
* INOUT : br_0_197 
* INOUT : bl_0_198 
* INOUT : br_0_198 
* INOUT : bl_0_199 
* INOUT : br_0_199 
* INOUT : bl_0_200 
* INOUT : br_0_200 
* INOUT : bl_0_201 
* INOUT : br_0_201 
* INOUT : bl_0_202 
* INOUT : br_0_202 
* INOUT : bl_0_203 
* INOUT : br_0_203 
* INOUT : bl_0_204 
* INOUT : br_0_204 
* INOUT : bl_0_205 
* INOUT : br_0_205 
* INOUT : bl_0_206 
* INOUT : br_0_206 
* INOUT : bl_0_207 
* INOUT : br_0_207 
* INOUT : bl_0_208 
* INOUT : br_0_208 
* INOUT : bl_0_209 
* INOUT : br_0_209 
* INOUT : bl_0_210 
* INOUT : br_0_210 
* INOUT : bl_0_211 
* INOUT : br_0_211 
* INOUT : bl_0_212 
* INOUT : br_0_212 
* INOUT : bl_0_213 
* INOUT : br_0_213 
* INOUT : bl_0_214 
* INOUT : br_0_214 
* INOUT : bl_0_215 
* INOUT : br_0_215 
* INOUT : bl_0_216 
* INOUT : br_0_216 
* INOUT : bl_0_217 
* INOUT : br_0_217 
* INOUT : bl_0_218 
* INOUT : br_0_218 
* INOUT : bl_0_219 
* INOUT : br_0_219 
* INOUT : bl_0_220 
* INOUT : br_0_220 
* INOUT : bl_0_221 
* INOUT : br_0_221 
* INOUT : bl_0_222 
* INOUT : br_0_222 
* INOUT : bl_0_223 
* INOUT : br_0_223 
* INOUT : bl_0_224 
* INOUT : br_0_224 
* INOUT : bl_0_225 
* INOUT : br_0_225 
* INOUT : bl_0_226 
* INOUT : br_0_226 
* INOUT : bl_0_227 
* INOUT : br_0_227 
* INOUT : bl_0_228 
* INOUT : br_0_228 
* INOUT : bl_0_229 
* INOUT : br_0_229 
* INOUT : bl_0_230 
* INOUT : br_0_230 
* INOUT : bl_0_231 
* INOUT : br_0_231 
* INOUT : bl_0_232 
* INOUT : br_0_232 
* INOUT : bl_0_233 
* INOUT : br_0_233 
* INOUT : bl_0_234 
* INOUT : br_0_234 
* INOUT : bl_0_235 
* INOUT : br_0_235 
* INOUT : bl_0_236 
* INOUT : br_0_236 
* INOUT : bl_0_237 
* INOUT : br_0_237 
* INOUT : bl_0_238 
* INOUT : br_0_238 
* INOUT : bl_0_239 
* INOUT : br_0_239 
* INOUT : bl_0_240 
* INOUT : br_0_240 
* INOUT : bl_0_241 
* INOUT : br_0_241 
* INOUT : bl_0_242 
* INOUT : br_0_242 
* INOUT : bl_0_243 
* INOUT : br_0_243 
* INOUT : bl_0_244 
* INOUT : br_0_244 
* INOUT : bl_0_245 
* INOUT : br_0_245 
* INOUT : bl_0_246 
* INOUT : br_0_246 
* INOUT : bl_0_247 
* INOUT : br_0_247 
* INOUT : bl_0_248 
* INOUT : br_0_248 
* INOUT : bl_0_249 
* INOUT : br_0_249 
* INOUT : bl_0_250 
* INOUT : br_0_250 
* INOUT : bl_0_251 
* INOUT : br_0_251 
* INOUT : bl_0_252 
* INOUT : br_0_252 
* INOUT : bl_0_253 
* INOUT : br_0_253 
* INOUT : bl_0_254 
* INOUT : br_0_254 
* INOUT : bl_0_255 
* INOUT : br_0_255 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* INPUT : wl_0_33 
* INPUT : wl_0_34 
* INPUT : wl_0_35 
* INPUT : wl_0_36 
* INPUT : wl_0_37 
* INPUT : wl_0_38 
* INPUT : wl_0_39 
* INPUT : wl_0_40 
* INPUT : wl_0_41 
* INPUT : wl_0_42 
* INPUT : wl_0_43 
* INPUT : wl_0_44 
* INPUT : wl_0_45 
* INPUT : wl_0_46 
* INPUT : wl_0_47 
* INPUT : wl_0_48 
* INPUT : wl_0_49 
* INPUT : wl_0_50 
* INPUT : wl_0_51 
* INPUT : wl_0_52 
* INPUT : wl_0_53 
* INPUT : wl_0_54 
* INPUT : wl_0_55 
* INPUT : wl_0_56 
* INPUT : wl_0_57 
* INPUT : wl_0_58 
* INPUT : wl_0_59 
* INPUT : wl_0_60 
* INPUT : wl_0_61 
* INPUT : wl_0_62 
* INPUT : wl_0_63 
* INPUT : wl_0_64 
* INPUT : wl_0_65 
* INPUT : wl_0_66 
* INPUT : wl_0_67 
* INPUT : wl_0_68 
* INPUT : wl_0_69 
* INPUT : wl_0_70 
* INPUT : wl_0_71 
* INPUT : wl_0_72 
* INPUT : wl_0_73 
* INPUT : wl_0_74 
* INPUT : wl_0_75 
* INPUT : wl_0_76 
* INPUT : wl_0_77 
* INPUT : wl_0_78 
* INPUT : wl_0_79 
* INPUT : wl_0_80 
* INPUT : wl_0_81 
* INPUT : wl_0_82 
* INPUT : wl_0_83 
* INPUT : wl_0_84 
* INPUT : wl_0_85 
* INPUT : wl_0_86 
* INPUT : wl_0_87 
* INPUT : wl_0_88 
* INPUT : wl_0_89 
* INPUT : wl_0_90 
* INPUT : wl_0_91 
* INPUT : wl_0_92 
* INPUT : wl_0_93 
* INPUT : wl_0_94 
* INPUT : wl_0_95 
* INPUT : wl_0_96 
* INPUT : wl_0_97 
* INPUT : wl_0_98 
* INPUT : wl_0_99 
* INPUT : wl_0_100 
* INPUT : wl_0_101 
* INPUT : wl_0_102 
* INPUT : wl_0_103 
* INPUT : wl_0_104 
* INPUT : wl_0_105 
* INPUT : wl_0_106 
* INPUT : wl_0_107 
* INPUT : wl_0_108 
* INPUT : wl_0_109 
* INPUT : wl_0_110 
* INPUT : wl_0_111 
* INPUT : wl_0_112 
* INPUT : wl_0_113 
* INPUT : wl_0_114 
* INPUT : wl_0_115 
* INPUT : wl_0_116 
* INPUT : wl_0_117 
* INPUT : wl_0_118 
* INPUT : wl_0_119 
* INPUT : wl_0_120 
* INPUT : wl_0_121 
* INPUT : wl_0_122 
* INPUT : wl_0_123 
* INPUT : wl_0_124 
* INPUT : wl_0_125 
* INPUT : wl_0_126 
* INPUT : wl_0_127 
* POWER : vdd 
* GROUND: gnd 
* rows: 128 cols: 256
Xbit_r0_c0
+ bl_0_0 br_0_0 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c0
+ bl_0_0 br_0_0 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c0
+ bl_0_0 br_0_0 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c0
+ bl_0_0 br_0_0 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c0
+ bl_0_0 br_0_0 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c0
+ bl_0_0 br_0_0 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c0
+ bl_0_0 br_0_0 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c0
+ bl_0_0 br_0_0 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c0
+ bl_0_0 br_0_0 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c0
+ bl_0_0 br_0_0 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c0
+ bl_0_0 br_0_0 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c0
+ bl_0_0 br_0_0 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c0
+ bl_0_0 br_0_0 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c0
+ bl_0_0 br_0_0 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c0
+ bl_0_0 br_0_0 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c0
+ bl_0_0 br_0_0 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c0
+ bl_0_0 br_0_0 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c0
+ bl_0_0 br_0_0 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c0
+ bl_0_0 br_0_0 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c0
+ bl_0_0 br_0_0 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c0
+ bl_0_0 br_0_0 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c0
+ bl_0_0 br_0_0 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c0
+ bl_0_0 br_0_0 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c0
+ bl_0_0 br_0_0 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c0
+ bl_0_0 br_0_0 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c0
+ bl_0_0 br_0_0 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c0
+ bl_0_0 br_0_0 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c0
+ bl_0_0 br_0_0 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c0
+ bl_0_0 br_0_0 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c0
+ bl_0_0 br_0_0 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c0
+ bl_0_0 br_0_0 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c0
+ bl_0_0 br_0_0 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c0
+ bl_0_0 br_0_0 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c0
+ bl_0_0 br_0_0 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c0
+ bl_0_0 br_0_0 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c0
+ bl_0_0 br_0_0 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c0
+ bl_0_0 br_0_0 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c0
+ bl_0_0 br_0_0 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c0
+ bl_0_0 br_0_0 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c0
+ bl_0_0 br_0_0 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c0
+ bl_0_0 br_0_0 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c0
+ bl_0_0 br_0_0 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c0
+ bl_0_0 br_0_0 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c0
+ bl_0_0 br_0_0 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c0
+ bl_0_0 br_0_0 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r45_c0
+ bl_0_0 br_0_0 wl_0_45 vdd gnd
+ cell_1rw
Xbit_r46_c0
+ bl_0_0 br_0_0 wl_0_46 vdd gnd
+ cell_1rw
Xbit_r47_c0
+ bl_0_0 br_0_0 wl_0_47 vdd gnd
+ cell_1rw
Xbit_r48_c0
+ bl_0_0 br_0_0 wl_0_48 vdd gnd
+ cell_1rw
Xbit_r49_c0
+ bl_0_0 br_0_0 wl_0_49 vdd gnd
+ cell_1rw
Xbit_r50_c0
+ bl_0_0 br_0_0 wl_0_50 vdd gnd
+ cell_1rw
Xbit_r51_c0
+ bl_0_0 br_0_0 wl_0_51 vdd gnd
+ cell_1rw
Xbit_r52_c0
+ bl_0_0 br_0_0 wl_0_52 vdd gnd
+ cell_1rw
Xbit_r53_c0
+ bl_0_0 br_0_0 wl_0_53 vdd gnd
+ cell_1rw
Xbit_r54_c0
+ bl_0_0 br_0_0 wl_0_54 vdd gnd
+ cell_1rw
Xbit_r55_c0
+ bl_0_0 br_0_0 wl_0_55 vdd gnd
+ cell_1rw
Xbit_r56_c0
+ bl_0_0 br_0_0 wl_0_56 vdd gnd
+ cell_1rw
Xbit_r57_c0
+ bl_0_0 br_0_0 wl_0_57 vdd gnd
+ cell_1rw
Xbit_r58_c0
+ bl_0_0 br_0_0 wl_0_58 vdd gnd
+ cell_1rw
Xbit_r59_c0
+ bl_0_0 br_0_0 wl_0_59 vdd gnd
+ cell_1rw
Xbit_r60_c0
+ bl_0_0 br_0_0 wl_0_60 vdd gnd
+ cell_1rw
Xbit_r61_c0
+ bl_0_0 br_0_0 wl_0_61 vdd gnd
+ cell_1rw
Xbit_r62_c0
+ bl_0_0 br_0_0 wl_0_62 vdd gnd
+ cell_1rw
Xbit_r63_c0
+ bl_0_0 br_0_0 wl_0_63 vdd gnd
+ cell_1rw
Xbit_r64_c0
+ bl_0_0 br_0_0 wl_0_64 vdd gnd
+ cell_1rw
Xbit_r65_c0
+ bl_0_0 br_0_0 wl_0_65 vdd gnd
+ cell_1rw
Xbit_r66_c0
+ bl_0_0 br_0_0 wl_0_66 vdd gnd
+ cell_1rw
Xbit_r67_c0
+ bl_0_0 br_0_0 wl_0_67 vdd gnd
+ cell_1rw
Xbit_r68_c0
+ bl_0_0 br_0_0 wl_0_68 vdd gnd
+ cell_1rw
Xbit_r69_c0
+ bl_0_0 br_0_0 wl_0_69 vdd gnd
+ cell_1rw
Xbit_r70_c0
+ bl_0_0 br_0_0 wl_0_70 vdd gnd
+ cell_1rw
Xbit_r71_c0
+ bl_0_0 br_0_0 wl_0_71 vdd gnd
+ cell_1rw
Xbit_r72_c0
+ bl_0_0 br_0_0 wl_0_72 vdd gnd
+ cell_1rw
Xbit_r73_c0
+ bl_0_0 br_0_0 wl_0_73 vdd gnd
+ cell_1rw
Xbit_r74_c0
+ bl_0_0 br_0_0 wl_0_74 vdd gnd
+ cell_1rw
Xbit_r75_c0
+ bl_0_0 br_0_0 wl_0_75 vdd gnd
+ cell_1rw
Xbit_r76_c0
+ bl_0_0 br_0_0 wl_0_76 vdd gnd
+ cell_1rw
Xbit_r77_c0
+ bl_0_0 br_0_0 wl_0_77 vdd gnd
+ cell_1rw
Xbit_r78_c0
+ bl_0_0 br_0_0 wl_0_78 vdd gnd
+ cell_1rw
Xbit_r79_c0
+ bl_0_0 br_0_0 wl_0_79 vdd gnd
+ cell_1rw
Xbit_r80_c0
+ bl_0_0 br_0_0 wl_0_80 vdd gnd
+ cell_1rw
Xbit_r81_c0
+ bl_0_0 br_0_0 wl_0_81 vdd gnd
+ cell_1rw
Xbit_r82_c0
+ bl_0_0 br_0_0 wl_0_82 vdd gnd
+ cell_1rw
Xbit_r83_c0
+ bl_0_0 br_0_0 wl_0_83 vdd gnd
+ cell_1rw
Xbit_r84_c0
+ bl_0_0 br_0_0 wl_0_84 vdd gnd
+ cell_1rw
Xbit_r85_c0
+ bl_0_0 br_0_0 wl_0_85 vdd gnd
+ cell_1rw
Xbit_r86_c0
+ bl_0_0 br_0_0 wl_0_86 vdd gnd
+ cell_1rw
Xbit_r87_c0
+ bl_0_0 br_0_0 wl_0_87 vdd gnd
+ cell_1rw
Xbit_r88_c0
+ bl_0_0 br_0_0 wl_0_88 vdd gnd
+ cell_1rw
Xbit_r89_c0
+ bl_0_0 br_0_0 wl_0_89 vdd gnd
+ cell_1rw
Xbit_r90_c0
+ bl_0_0 br_0_0 wl_0_90 vdd gnd
+ cell_1rw
Xbit_r91_c0
+ bl_0_0 br_0_0 wl_0_91 vdd gnd
+ cell_1rw
Xbit_r92_c0
+ bl_0_0 br_0_0 wl_0_92 vdd gnd
+ cell_1rw
Xbit_r93_c0
+ bl_0_0 br_0_0 wl_0_93 vdd gnd
+ cell_1rw
Xbit_r94_c0
+ bl_0_0 br_0_0 wl_0_94 vdd gnd
+ cell_1rw
Xbit_r95_c0
+ bl_0_0 br_0_0 wl_0_95 vdd gnd
+ cell_1rw
Xbit_r96_c0
+ bl_0_0 br_0_0 wl_0_96 vdd gnd
+ cell_1rw
Xbit_r97_c0
+ bl_0_0 br_0_0 wl_0_97 vdd gnd
+ cell_1rw
Xbit_r98_c0
+ bl_0_0 br_0_0 wl_0_98 vdd gnd
+ cell_1rw
Xbit_r99_c0
+ bl_0_0 br_0_0 wl_0_99 vdd gnd
+ cell_1rw
Xbit_r100_c0
+ bl_0_0 br_0_0 wl_0_100 vdd gnd
+ cell_1rw
Xbit_r101_c0
+ bl_0_0 br_0_0 wl_0_101 vdd gnd
+ cell_1rw
Xbit_r102_c0
+ bl_0_0 br_0_0 wl_0_102 vdd gnd
+ cell_1rw
Xbit_r103_c0
+ bl_0_0 br_0_0 wl_0_103 vdd gnd
+ cell_1rw
Xbit_r104_c0
+ bl_0_0 br_0_0 wl_0_104 vdd gnd
+ cell_1rw
Xbit_r105_c0
+ bl_0_0 br_0_0 wl_0_105 vdd gnd
+ cell_1rw
Xbit_r106_c0
+ bl_0_0 br_0_0 wl_0_106 vdd gnd
+ cell_1rw
Xbit_r107_c0
+ bl_0_0 br_0_0 wl_0_107 vdd gnd
+ cell_1rw
Xbit_r108_c0
+ bl_0_0 br_0_0 wl_0_108 vdd gnd
+ cell_1rw
Xbit_r109_c0
+ bl_0_0 br_0_0 wl_0_109 vdd gnd
+ cell_1rw
Xbit_r110_c0
+ bl_0_0 br_0_0 wl_0_110 vdd gnd
+ cell_1rw
Xbit_r111_c0
+ bl_0_0 br_0_0 wl_0_111 vdd gnd
+ cell_1rw
Xbit_r112_c0
+ bl_0_0 br_0_0 wl_0_112 vdd gnd
+ cell_1rw
Xbit_r113_c0
+ bl_0_0 br_0_0 wl_0_113 vdd gnd
+ cell_1rw
Xbit_r114_c0
+ bl_0_0 br_0_0 wl_0_114 vdd gnd
+ cell_1rw
Xbit_r115_c0
+ bl_0_0 br_0_0 wl_0_115 vdd gnd
+ cell_1rw
Xbit_r116_c0
+ bl_0_0 br_0_0 wl_0_116 vdd gnd
+ cell_1rw
Xbit_r117_c0
+ bl_0_0 br_0_0 wl_0_117 vdd gnd
+ cell_1rw
Xbit_r118_c0
+ bl_0_0 br_0_0 wl_0_118 vdd gnd
+ cell_1rw
Xbit_r119_c0
+ bl_0_0 br_0_0 wl_0_119 vdd gnd
+ cell_1rw
Xbit_r120_c0
+ bl_0_0 br_0_0 wl_0_120 vdd gnd
+ cell_1rw
Xbit_r121_c0
+ bl_0_0 br_0_0 wl_0_121 vdd gnd
+ cell_1rw
Xbit_r122_c0
+ bl_0_0 br_0_0 wl_0_122 vdd gnd
+ cell_1rw
Xbit_r123_c0
+ bl_0_0 br_0_0 wl_0_123 vdd gnd
+ cell_1rw
Xbit_r124_c0
+ bl_0_0 br_0_0 wl_0_124 vdd gnd
+ cell_1rw
Xbit_r125_c0
+ bl_0_0 br_0_0 wl_0_125 vdd gnd
+ cell_1rw
Xbit_r126_c0
+ bl_0_0 br_0_0 wl_0_126 vdd gnd
+ cell_1rw
Xbit_r127_c0
+ bl_0_0 br_0_0 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c1
+ bl_0_1 br_0_1 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c1
*+ bl_0_1 br_0_1 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c1
*+ bl_0_1 br_0_1 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c1
*+ bl_0_1 br_0_1 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c1
*+ bl_0_1 br_0_1 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c1
*+ bl_0_1 br_0_1 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c1
*+ bl_0_1 br_0_1 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c1
*+ bl_0_1 br_0_1 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c1
*+ bl_0_1 br_0_1 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c1
*+ bl_0_1 br_0_1 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c1
*+ bl_0_1 br_0_1 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c1
*+ bl_0_1 br_0_1 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c1
*+ bl_0_1 br_0_1 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c1
*+ bl_0_1 br_0_1 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c1
*+ bl_0_1 br_0_1 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c1
*+ bl_0_1 br_0_1 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c1
*+ bl_0_1 br_0_1 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c1
*+ bl_0_1 br_0_1 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c1
*+ bl_0_1 br_0_1 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c1
*+ bl_0_1 br_0_1 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c1
*+ bl_0_1 br_0_1 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c1
*+ bl_0_1 br_0_1 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c1
*+ bl_0_1 br_0_1 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c1
*+ bl_0_1 br_0_1 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c1
*+ bl_0_1 br_0_1 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c1
*+ bl_0_1 br_0_1 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c1
*+ bl_0_1 br_0_1 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c1
*+ bl_0_1 br_0_1 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c1
*+ bl_0_1 br_0_1 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c1
*+ bl_0_1 br_0_1 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c1
*+ bl_0_1 br_0_1 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c1
*+ bl_0_1 br_0_1 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c1
*+ bl_0_1 br_0_1 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c1
*+ bl_0_1 br_0_1 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c1
*+ bl_0_1 br_0_1 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c1
*+ bl_0_1 br_0_1 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c1
*+ bl_0_1 br_0_1 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c1
*+ bl_0_1 br_0_1 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c1
*+ bl_0_1 br_0_1 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c1
*+ bl_0_1 br_0_1 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c1
*+ bl_0_1 br_0_1 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c1
*+ bl_0_1 br_0_1 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c1
*+ bl_0_1 br_0_1 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c1
*+ bl_0_1 br_0_1 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c1
*+ bl_0_1 br_0_1 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c1
*+ bl_0_1 br_0_1 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c1
*+ bl_0_1 br_0_1 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c1
*+ bl_0_1 br_0_1 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c1
*+ bl_0_1 br_0_1 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c1
*+ bl_0_1 br_0_1 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c1
*+ bl_0_1 br_0_1 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c1
*+ bl_0_1 br_0_1 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c1
*+ bl_0_1 br_0_1 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c1
*+ bl_0_1 br_0_1 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c1
*+ bl_0_1 br_0_1 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c1
*+ bl_0_1 br_0_1 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c1
*+ bl_0_1 br_0_1 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c1
*+ bl_0_1 br_0_1 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c1
*+ bl_0_1 br_0_1 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c1
*+ bl_0_1 br_0_1 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c1
*+ bl_0_1 br_0_1 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c1
*+ bl_0_1 br_0_1 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c1
*+ bl_0_1 br_0_1 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c1
*+ bl_0_1 br_0_1 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c1
*+ bl_0_1 br_0_1 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c1
*+ bl_0_1 br_0_1 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c1
*+ bl_0_1 br_0_1 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c1
*+ bl_0_1 br_0_1 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c1
*+ bl_0_1 br_0_1 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c1
*+ bl_0_1 br_0_1 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c1
*+ bl_0_1 br_0_1 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c1
*+ bl_0_1 br_0_1 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c1
*+ bl_0_1 br_0_1 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c1
*+ bl_0_1 br_0_1 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c1
*+ bl_0_1 br_0_1 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c1
*+ bl_0_1 br_0_1 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c1
*+ bl_0_1 br_0_1 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c1
*+ bl_0_1 br_0_1 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c1
*+ bl_0_1 br_0_1 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c1
*+ bl_0_1 br_0_1 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c1
*+ bl_0_1 br_0_1 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c1
*+ bl_0_1 br_0_1 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c1
*+ bl_0_1 br_0_1 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c1
*+ bl_0_1 br_0_1 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c1
*+ bl_0_1 br_0_1 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c1
*+ bl_0_1 br_0_1 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c1
*+ bl_0_1 br_0_1 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c1
*+ bl_0_1 br_0_1 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c1
*+ bl_0_1 br_0_1 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c1
*+ bl_0_1 br_0_1 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c1
*+ bl_0_1 br_0_1 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c1
*+ bl_0_1 br_0_1 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c1
*+ bl_0_1 br_0_1 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c1
*+ bl_0_1 br_0_1 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c1
*+ bl_0_1 br_0_1 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c1
*+ bl_0_1 br_0_1 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c1
*+ bl_0_1 br_0_1 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c1
*+ bl_0_1 br_0_1 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c1
*+ bl_0_1 br_0_1 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c1
*+ bl_0_1 br_0_1 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c1
*+ bl_0_1 br_0_1 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c1
*+ bl_0_1 br_0_1 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c1
*+ bl_0_1 br_0_1 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c1
*+ bl_0_1 br_0_1 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c1
*+ bl_0_1 br_0_1 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c1
*+ bl_0_1 br_0_1 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c1
*+ bl_0_1 br_0_1 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c1
*+ bl_0_1 br_0_1 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c1
*+ bl_0_1 br_0_1 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c1
*+ bl_0_1 br_0_1 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c1
*+ bl_0_1 br_0_1 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c1
*+ bl_0_1 br_0_1 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c1
*+ bl_0_1 br_0_1 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c1
*+ bl_0_1 br_0_1 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c1
*+ bl_0_1 br_0_1 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c1
*+ bl_0_1 br_0_1 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c1
*+ bl_0_1 br_0_1 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c1
*+ bl_0_1 br_0_1 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c1
*+ bl_0_1 br_0_1 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c1
*+ bl_0_1 br_0_1 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c1
*+ bl_0_1 br_0_1 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c1
*+ bl_0_1 br_0_1 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c1
*+ bl_0_1 br_0_1 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c1
*+ bl_0_1 br_0_1 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c1
*+ bl_0_1 br_0_1 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c1
*+ bl_0_1 br_0_1 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c1
*+ bl_0_1 br_0_1 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c1
+ bl_0_1 br_0_1 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c2
+ bl_0_2 br_0_2 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c2
*+ bl_0_2 br_0_2 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c2
*+ bl_0_2 br_0_2 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c2
*+ bl_0_2 br_0_2 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c2
*+ bl_0_2 br_0_2 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c2
*+ bl_0_2 br_0_2 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c2
*+ bl_0_2 br_0_2 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c2
*+ bl_0_2 br_0_2 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c2
*+ bl_0_2 br_0_2 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c2
*+ bl_0_2 br_0_2 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c2
*+ bl_0_2 br_0_2 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c2
*+ bl_0_2 br_0_2 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c2
*+ bl_0_2 br_0_2 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c2
*+ bl_0_2 br_0_2 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c2
*+ bl_0_2 br_0_2 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c2
*+ bl_0_2 br_0_2 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c2
*+ bl_0_2 br_0_2 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c2
*+ bl_0_2 br_0_2 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c2
*+ bl_0_2 br_0_2 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c2
*+ bl_0_2 br_0_2 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c2
*+ bl_0_2 br_0_2 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c2
*+ bl_0_2 br_0_2 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c2
*+ bl_0_2 br_0_2 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c2
*+ bl_0_2 br_0_2 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c2
*+ bl_0_2 br_0_2 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c2
*+ bl_0_2 br_0_2 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c2
*+ bl_0_2 br_0_2 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c2
*+ bl_0_2 br_0_2 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c2
*+ bl_0_2 br_0_2 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c2
*+ bl_0_2 br_0_2 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c2
*+ bl_0_2 br_0_2 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c2
*+ bl_0_2 br_0_2 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c2
*+ bl_0_2 br_0_2 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c2
*+ bl_0_2 br_0_2 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c2
*+ bl_0_2 br_0_2 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c2
*+ bl_0_2 br_0_2 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c2
*+ bl_0_2 br_0_2 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c2
*+ bl_0_2 br_0_2 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c2
*+ bl_0_2 br_0_2 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c2
*+ bl_0_2 br_0_2 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c2
*+ bl_0_2 br_0_2 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c2
*+ bl_0_2 br_0_2 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c2
*+ bl_0_2 br_0_2 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c2
*+ bl_0_2 br_0_2 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c2
*+ bl_0_2 br_0_2 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c2
*+ bl_0_2 br_0_2 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c2
*+ bl_0_2 br_0_2 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c2
*+ bl_0_2 br_0_2 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c2
*+ bl_0_2 br_0_2 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c2
*+ bl_0_2 br_0_2 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c2
*+ bl_0_2 br_0_2 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c2
*+ bl_0_2 br_0_2 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c2
*+ bl_0_2 br_0_2 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c2
*+ bl_0_2 br_0_2 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c2
*+ bl_0_2 br_0_2 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c2
*+ bl_0_2 br_0_2 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c2
*+ bl_0_2 br_0_2 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c2
*+ bl_0_2 br_0_2 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c2
*+ bl_0_2 br_0_2 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c2
*+ bl_0_2 br_0_2 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c2
*+ bl_0_2 br_0_2 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c2
*+ bl_0_2 br_0_2 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c2
*+ bl_0_2 br_0_2 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c2
*+ bl_0_2 br_0_2 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c2
*+ bl_0_2 br_0_2 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c2
*+ bl_0_2 br_0_2 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c2
*+ bl_0_2 br_0_2 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c2
*+ bl_0_2 br_0_2 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c2
*+ bl_0_2 br_0_2 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c2
*+ bl_0_2 br_0_2 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c2
*+ bl_0_2 br_0_2 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c2
*+ bl_0_2 br_0_2 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c2
*+ bl_0_2 br_0_2 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c2
*+ bl_0_2 br_0_2 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c2
*+ bl_0_2 br_0_2 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c2
*+ bl_0_2 br_0_2 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c2
*+ bl_0_2 br_0_2 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c2
*+ bl_0_2 br_0_2 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c2
*+ bl_0_2 br_0_2 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c2
*+ bl_0_2 br_0_2 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c2
*+ bl_0_2 br_0_2 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c2
*+ bl_0_2 br_0_2 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c2
*+ bl_0_2 br_0_2 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c2
*+ bl_0_2 br_0_2 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c2
*+ bl_0_2 br_0_2 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c2
*+ bl_0_2 br_0_2 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c2
*+ bl_0_2 br_0_2 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c2
*+ bl_0_2 br_0_2 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c2
*+ bl_0_2 br_0_2 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c2
*+ bl_0_2 br_0_2 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c2
*+ bl_0_2 br_0_2 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c2
*+ bl_0_2 br_0_2 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c2
*+ bl_0_2 br_0_2 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c2
*+ bl_0_2 br_0_2 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c2
*+ bl_0_2 br_0_2 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c2
*+ bl_0_2 br_0_2 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c2
*+ bl_0_2 br_0_2 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c2
*+ bl_0_2 br_0_2 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c2
*+ bl_0_2 br_0_2 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c2
*+ bl_0_2 br_0_2 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c2
*+ bl_0_2 br_0_2 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c2
*+ bl_0_2 br_0_2 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c2
*+ bl_0_2 br_0_2 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c2
*+ bl_0_2 br_0_2 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c2
*+ bl_0_2 br_0_2 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c2
*+ bl_0_2 br_0_2 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c2
*+ bl_0_2 br_0_2 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c2
*+ bl_0_2 br_0_2 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c2
*+ bl_0_2 br_0_2 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c2
*+ bl_0_2 br_0_2 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c2
*+ bl_0_2 br_0_2 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c2
*+ bl_0_2 br_0_2 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c2
*+ bl_0_2 br_0_2 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c2
*+ bl_0_2 br_0_2 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c2
*+ bl_0_2 br_0_2 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c2
*+ bl_0_2 br_0_2 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c2
*+ bl_0_2 br_0_2 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c2
*+ bl_0_2 br_0_2 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c2
*+ bl_0_2 br_0_2 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c2
*+ bl_0_2 br_0_2 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c2
*+ bl_0_2 br_0_2 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c2
*+ bl_0_2 br_0_2 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c2
*+ bl_0_2 br_0_2 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c2
*+ bl_0_2 br_0_2 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c2
*+ bl_0_2 br_0_2 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c2
*+ bl_0_2 br_0_2 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c2
*+ bl_0_2 br_0_2 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c2
+ bl_0_2 br_0_2 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c3
+ bl_0_3 br_0_3 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c3
*+ bl_0_3 br_0_3 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c3
*+ bl_0_3 br_0_3 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c3
*+ bl_0_3 br_0_3 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c3
*+ bl_0_3 br_0_3 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c3
*+ bl_0_3 br_0_3 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c3
*+ bl_0_3 br_0_3 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c3
*+ bl_0_3 br_0_3 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c3
*+ bl_0_3 br_0_3 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c3
*+ bl_0_3 br_0_3 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c3
*+ bl_0_3 br_0_3 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c3
*+ bl_0_3 br_0_3 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c3
*+ bl_0_3 br_0_3 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c3
*+ bl_0_3 br_0_3 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c3
*+ bl_0_3 br_0_3 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c3
*+ bl_0_3 br_0_3 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c3
*+ bl_0_3 br_0_3 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c3
*+ bl_0_3 br_0_3 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c3
*+ bl_0_3 br_0_3 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c3
*+ bl_0_3 br_0_3 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c3
*+ bl_0_3 br_0_3 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c3
*+ bl_0_3 br_0_3 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c3
*+ bl_0_3 br_0_3 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c3
*+ bl_0_3 br_0_3 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c3
*+ bl_0_3 br_0_3 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c3
*+ bl_0_3 br_0_3 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c3
*+ bl_0_3 br_0_3 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c3
*+ bl_0_3 br_0_3 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c3
*+ bl_0_3 br_0_3 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c3
*+ bl_0_3 br_0_3 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c3
*+ bl_0_3 br_0_3 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c3
*+ bl_0_3 br_0_3 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c3
*+ bl_0_3 br_0_3 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c3
*+ bl_0_3 br_0_3 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c3
*+ bl_0_3 br_0_3 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c3
*+ bl_0_3 br_0_3 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c3
*+ bl_0_3 br_0_3 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c3
*+ bl_0_3 br_0_3 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c3
*+ bl_0_3 br_0_3 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c3
*+ bl_0_3 br_0_3 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c3
*+ bl_0_3 br_0_3 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c3
*+ bl_0_3 br_0_3 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c3
*+ bl_0_3 br_0_3 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c3
*+ bl_0_3 br_0_3 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c3
*+ bl_0_3 br_0_3 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c3
*+ bl_0_3 br_0_3 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c3
*+ bl_0_3 br_0_3 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c3
*+ bl_0_3 br_0_3 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c3
*+ bl_0_3 br_0_3 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c3
*+ bl_0_3 br_0_3 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c3
*+ bl_0_3 br_0_3 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c3
*+ bl_0_3 br_0_3 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c3
*+ bl_0_3 br_0_3 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c3
*+ bl_0_3 br_0_3 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c3
*+ bl_0_3 br_0_3 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c3
*+ bl_0_3 br_0_3 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c3
*+ bl_0_3 br_0_3 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c3
*+ bl_0_3 br_0_3 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c3
*+ bl_0_3 br_0_3 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c3
*+ bl_0_3 br_0_3 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c3
*+ bl_0_3 br_0_3 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c3
*+ bl_0_3 br_0_3 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c3
*+ bl_0_3 br_0_3 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c3
*+ bl_0_3 br_0_3 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c3
*+ bl_0_3 br_0_3 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c3
*+ bl_0_3 br_0_3 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c3
*+ bl_0_3 br_0_3 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c3
*+ bl_0_3 br_0_3 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c3
*+ bl_0_3 br_0_3 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c3
*+ bl_0_3 br_0_3 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c3
*+ bl_0_3 br_0_3 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c3
*+ bl_0_3 br_0_3 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c3
*+ bl_0_3 br_0_3 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c3
*+ bl_0_3 br_0_3 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c3
*+ bl_0_3 br_0_3 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c3
*+ bl_0_3 br_0_3 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c3
*+ bl_0_3 br_0_3 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c3
*+ bl_0_3 br_0_3 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c3
*+ bl_0_3 br_0_3 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c3
*+ bl_0_3 br_0_3 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c3
*+ bl_0_3 br_0_3 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c3
*+ bl_0_3 br_0_3 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c3
*+ bl_0_3 br_0_3 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c3
*+ bl_0_3 br_0_3 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c3
*+ bl_0_3 br_0_3 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c3
*+ bl_0_3 br_0_3 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c3
*+ bl_0_3 br_0_3 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c3
*+ bl_0_3 br_0_3 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c3
*+ bl_0_3 br_0_3 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c3
*+ bl_0_3 br_0_3 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c3
*+ bl_0_3 br_0_3 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c3
*+ bl_0_3 br_0_3 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c3
*+ bl_0_3 br_0_3 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c3
*+ bl_0_3 br_0_3 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c3
*+ bl_0_3 br_0_3 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c3
*+ bl_0_3 br_0_3 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c3
*+ bl_0_3 br_0_3 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c3
*+ bl_0_3 br_0_3 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c3
*+ bl_0_3 br_0_3 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c3
*+ bl_0_3 br_0_3 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c3
*+ bl_0_3 br_0_3 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c3
*+ bl_0_3 br_0_3 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c3
*+ bl_0_3 br_0_3 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c3
*+ bl_0_3 br_0_3 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c3
*+ bl_0_3 br_0_3 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c3
*+ bl_0_3 br_0_3 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c3
*+ bl_0_3 br_0_3 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c3
*+ bl_0_3 br_0_3 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c3
*+ bl_0_3 br_0_3 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c3
*+ bl_0_3 br_0_3 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c3
*+ bl_0_3 br_0_3 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c3
*+ bl_0_3 br_0_3 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c3
*+ bl_0_3 br_0_3 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c3
*+ bl_0_3 br_0_3 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c3
*+ bl_0_3 br_0_3 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c3
*+ bl_0_3 br_0_3 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c3
*+ bl_0_3 br_0_3 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c3
*+ bl_0_3 br_0_3 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c3
*+ bl_0_3 br_0_3 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c3
*+ bl_0_3 br_0_3 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c3
*+ bl_0_3 br_0_3 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c3
*+ bl_0_3 br_0_3 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c3
*+ bl_0_3 br_0_3 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c3
*+ bl_0_3 br_0_3 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c3
*+ bl_0_3 br_0_3 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c3
*+ bl_0_3 br_0_3 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c3
*+ bl_0_3 br_0_3 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c3
+ bl_0_3 br_0_3 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c4
+ bl_0_4 br_0_4 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c4
*+ bl_0_4 br_0_4 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c4
*+ bl_0_4 br_0_4 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c4
*+ bl_0_4 br_0_4 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c4
*+ bl_0_4 br_0_4 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c4
*+ bl_0_4 br_0_4 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c4
*+ bl_0_4 br_0_4 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c4
*+ bl_0_4 br_0_4 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c4
*+ bl_0_4 br_0_4 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c4
*+ bl_0_4 br_0_4 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c4
*+ bl_0_4 br_0_4 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c4
*+ bl_0_4 br_0_4 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c4
*+ bl_0_4 br_0_4 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c4
*+ bl_0_4 br_0_4 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c4
*+ bl_0_4 br_0_4 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c4
*+ bl_0_4 br_0_4 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c4
*+ bl_0_4 br_0_4 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c4
*+ bl_0_4 br_0_4 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c4
*+ bl_0_4 br_0_4 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c4
*+ bl_0_4 br_0_4 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c4
*+ bl_0_4 br_0_4 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c4
*+ bl_0_4 br_0_4 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c4
*+ bl_0_4 br_0_4 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c4
*+ bl_0_4 br_0_4 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c4
*+ bl_0_4 br_0_4 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c4
*+ bl_0_4 br_0_4 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c4
*+ bl_0_4 br_0_4 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c4
*+ bl_0_4 br_0_4 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c4
*+ bl_0_4 br_0_4 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c4
*+ bl_0_4 br_0_4 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c4
*+ bl_0_4 br_0_4 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c4
*+ bl_0_4 br_0_4 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c4
*+ bl_0_4 br_0_4 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c4
*+ bl_0_4 br_0_4 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c4
*+ bl_0_4 br_0_4 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c4
*+ bl_0_4 br_0_4 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c4
*+ bl_0_4 br_0_4 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c4
*+ bl_0_4 br_0_4 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c4
*+ bl_0_4 br_0_4 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c4
*+ bl_0_4 br_0_4 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c4
*+ bl_0_4 br_0_4 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c4
*+ bl_0_4 br_0_4 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c4
*+ bl_0_4 br_0_4 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c4
*+ bl_0_4 br_0_4 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c4
*+ bl_0_4 br_0_4 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c4
*+ bl_0_4 br_0_4 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c4
*+ bl_0_4 br_0_4 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c4
*+ bl_0_4 br_0_4 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c4
*+ bl_0_4 br_0_4 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c4
*+ bl_0_4 br_0_4 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c4
*+ bl_0_4 br_0_4 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c4
*+ bl_0_4 br_0_4 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c4
*+ bl_0_4 br_0_4 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c4
*+ bl_0_4 br_0_4 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c4
*+ bl_0_4 br_0_4 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c4
*+ bl_0_4 br_0_4 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c4
*+ bl_0_4 br_0_4 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c4
*+ bl_0_4 br_0_4 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c4
*+ bl_0_4 br_0_4 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c4
*+ bl_0_4 br_0_4 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c4
*+ bl_0_4 br_0_4 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c4
*+ bl_0_4 br_0_4 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c4
*+ bl_0_4 br_0_4 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c4
*+ bl_0_4 br_0_4 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c4
*+ bl_0_4 br_0_4 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c4
*+ bl_0_4 br_0_4 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c4
*+ bl_0_4 br_0_4 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c4
*+ bl_0_4 br_0_4 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c4
*+ bl_0_4 br_0_4 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c4
*+ bl_0_4 br_0_4 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c4
*+ bl_0_4 br_0_4 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c4
*+ bl_0_4 br_0_4 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c4
*+ bl_0_4 br_0_4 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c4
*+ bl_0_4 br_0_4 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c4
*+ bl_0_4 br_0_4 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c4
*+ bl_0_4 br_0_4 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c4
*+ bl_0_4 br_0_4 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c4
*+ bl_0_4 br_0_4 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c4
*+ bl_0_4 br_0_4 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c4
*+ bl_0_4 br_0_4 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c4
*+ bl_0_4 br_0_4 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c4
*+ bl_0_4 br_0_4 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c4
*+ bl_0_4 br_0_4 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c4
*+ bl_0_4 br_0_4 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c4
*+ bl_0_4 br_0_4 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c4
*+ bl_0_4 br_0_4 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c4
*+ bl_0_4 br_0_4 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c4
*+ bl_0_4 br_0_4 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c4
*+ bl_0_4 br_0_4 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c4
*+ bl_0_4 br_0_4 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c4
*+ bl_0_4 br_0_4 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c4
*+ bl_0_4 br_0_4 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c4
*+ bl_0_4 br_0_4 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c4
*+ bl_0_4 br_0_4 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c4
*+ bl_0_4 br_0_4 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c4
*+ bl_0_4 br_0_4 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c4
*+ bl_0_4 br_0_4 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c4
*+ bl_0_4 br_0_4 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c4
*+ bl_0_4 br_0_4 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c4
*+ bl_0_4 br_0_4 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c4
*+ bl_0_4 br_0_4 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c4
*+ bl_0_4 br_0_4 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c4
*+ bl_0_4 br_0_4 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c4
*+ bl_0_4 br_0_4 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c4
*+ bl_0_4 br_0_4 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c4
*+ bl_0_4 br_0_4 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c4
*+ bl_0_4 br_0_4 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c4
*+ bl_0_4 br_0_4 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c4
*+ bl_0_4 br_0_4 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c4
*+ bl_0_4 br_0_4 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c4
*+ bl_0_4 br_0_4 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c4
*+ bl_0_4 br_0_4 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c4
*+ bl_0_4 br_0_4 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c4
*+ bl_0_4 br_0_4 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c4
*+ bl_0_4 br_0_4 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c4
*+ bl_0_4 br_0_4 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c4
*+ bl_0_4 br_0_4 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c4
*+ bl_0_4 br_0_4 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c4
*+ bl_0_4 br_0_4 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c4
*+ bl_0_4 br_0_4 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c4
*+ bl_0_4 br_0_4 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c4
*+ bl_0_4 br_0_4 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c4
*+ bl_0_4 br_0_4 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c4
*+ bl_0_4 br_0_4 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c4
*+ bl_0_4 br_0_4 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c4
*+ bl_0_4 br_0_4 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c4
*+ bl_0_4 br_0_4 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c4
+ bl_0_4 br_0_4 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c5
+ bl_0_5 br_0_5 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c5
*+ bl_0_5 br_0_5 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c5
*+ bl_0_5 br_0_5 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c5
*+ bl_0_5 br_0_5 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c5
*+ bl_0_5 br_0_5 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c5
*+ bl_0_5 br_0_5 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c5
*+ bl_0_5 br_0_5 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c5
*+ bl_0_5 br_0_5 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c5
*+ bl_0_5 br_0_5 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c5
*+ bl_0_5 br_0_5 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c5
*+ bl_0_5 br_0_5 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c5
*+ bl_0_5 br_0_5 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c5
*+ bl_0_5 br_0_5 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c5
*+ bl_0_5 br_0_5 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c5
*+ bl_0_5 br_0_5 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c5
*+ bl_0_5 br_0_5 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c5
*+ bl_0_5 br_0_5 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c5
*+ bl_0_5 br_0_5 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c5
*+ bl_0_5 br_0_5 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c5
*+ bl_0_5 br_0_5 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c5
*+ bl_0_5 br_0_5 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c5
*+ bl_0_5 br_0_5 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c5
*+ bl_0_5 br_0_5 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c5
*+ bl_0_5 br_0_5 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c5
*+ bl_0_5 br_0_5 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c5
*+ bl_0_5 br_0_5 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c5
*+ bl_0_5 br_0_5 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c5
*+ bl_0_5 br_0_5 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c5
*+ bl_0_5 br_0_5 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c5
*+ bl_0_5 br_0_5 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c5
*+ bl_0_5 br_0_5 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c5
*+ bl_0_5 br_0_5 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c5
*+ bl_0_5 br_0_5 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c5
*+ bl_0_5 br_0_5 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c5
*+ bl_0_5 br_0_5 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c5
*+ bl_0_5 br_0_5 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c5
*+ bl_0_5 br_0_5 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c5
*+ bl_0_5 br_0_5 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c5
*+ bl_0_5 br_0_5 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c5
*+ bl_0_5 br_0_5 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c5
*+ bl_0_5 br_0_5 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c5
*+ bl_0_5 br_0_5 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c5
*+ bl_0_5 br_0_5 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c5
*+ bl_0_5 br_0_5 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c5
*+ bl_0_5 br_0_5 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c5
*+ bl_0_5 br_0_5 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c5
*+ bl_0_5 br_0_5 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c5
*+ bl_0_5 br_0_5 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c5
*+ bl_0_5 br_0_5 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c5
*+ bl_0_5 br_0_5 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c5
*+ bl_0_5 br_0_5 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c5
*+ bl_0_5 br_0_5 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c5
*+ bl_0_5 br_0_5 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c5
*+ bl_0_5 br_0_5 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c5
*+ bl_0_5 br_0_5 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c5
*+ bl_0_5 br_0_5 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c5
*+ bl_0_5 br_0_5 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c5
*+ bl_0_5 br_0_5 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c5
*+ bl_0_5 br_0_5 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c5
*+ bl_0_5 br_0_5 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c5
*+ bl_0_5 br_0_5 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c5
*+ bl_0_5 br_0_5 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c5
*+ bl_0_5 br_0_5 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c5
*+ bl_0_5 br_0_5 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c5
*+ bl_0_5 br_0_5 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c5
*+ bl_0_5 br_0_5 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c5
*+ bl_0_5 br_0_5 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c5
*+ bl_0_5 br_0_5 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c5
*+ bl_0_5 br_0_5 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c5
*+ bl_0_5 br_0_5 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c5
*+ bl_0_5 br_0_5 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c5
*+ bl_0_5 br_0_5 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c5
*+ bl_0_5 br_0_5 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c5
*+ bl_0_5 br_0_5 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c5
*+ bl_0_5 br_0_5 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c5
*+ bl_0_5 br_0_5 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c5
*+ bl_0_5 br_0_5 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c5
*+ bl_0_5 br_0_5 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c5
*+ bl_0_5 br_0_5 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c5
*+ bl_0_5 br_0_5 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c5
*+ bl_0_5 br_0_5 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c5
*+ bl_0_5 br_0_5 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c5
*+ bl_0_5 br_0_5 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c5
*+ bl_0_5 br_0_5 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c5
*+ bl_0_5 br_0_5 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c5
*+ bl_0_5 br_0_5 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c5
*+ bl_0_5 br_0_5 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c5
*+ bl_0_5 br_0_5 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c5
*+ bl_0_5 br_0_5 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c5
*+ bl_0_5 br_0_5 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c5
*+ bl_0_5 br_0_5 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c5
*+ bl_0_5 br_0_5 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c5
*+ bl_0_5 br_0_5 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c5
*+ bl_0_5 br_0_5 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c5
*+ bl_0_5 br_0_5 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c5
*+ bl_0_5 br_0_5 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c5
*+ bl_0_5 br_0_5 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c5
*+ bl_0_5 br_0_5 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c5
*+ bl_0_5 br_0_5 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c5
*+ bl_0_5 br_0_5 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c5
*+ bl_0_5 br_0_5 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c5
*+ bl_0_5 br_0_5 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c5
*+ bl_0_5 br_0_5 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c5
*+ bl_0_5 br_0_5 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c5
*+ bl_0_5 br_0_5 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c5
*+ bl_0_5 br_0_5 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c5
*+ bl_0_5 br_0_5 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c5
*+ bl_0_5 br_0_5 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c5
*+ bl_0_5 br_0_5 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c5
*+ bl_0_5 br_0_5 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c5
*+ bl_0_5 br_0_5 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c5
*+ bl_0_5 br_0_5 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c5
*+ bl_0_5 br_0_5 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c5
*+ bl_0_5 br_0_5 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c5
*+ bl_0_5 br_0_5 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c5
*+ bl_0_5 br_0_5 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c5
*+ bl_0_5 br_0_5 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c5
*+ bl_0_5 br_0_5 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c5
*+ bl_0_5 br_0_5 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c5
*+ bl_0_5 br_0_5 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c5
*+ bl_0_5 br_0_5 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c5
*+ bl_0_5 br_0_5 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c5
*+ bl_0_5 br_0_5 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c5
*+ bl_0_5 br_0_5 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c5
*+ bl_0_5 br_0_5 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c5
*+ bl_0_5 br_0_5 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c5
*+ bl_0_5 br_0_5 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c5
+ bl_0_5 br_0_5 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c6
+ bl_0_6 br_0_6 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c6
*+ bl_0_6 br_0_6 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c6
*+ bl_0_6 br_0_6 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c6
*+ bl_0_6 br_0_6 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c6
*+ bl_0_6 br_0_6 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c6
*+ bl_0_6 br_0_6 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c6
*+ bl_0_6 br_0_6 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c6
*+ bl_0_6 br_0_6 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c6
*+ bl_0_6 br_0_6 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c6
*+ bl_0_6 br_0_6 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c6
*+ bl_0_6 br_0_6 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c6
*+ bl_0_6 br_0_6 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c6
*+ bl_0_6 br_0_6 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c6
*+ bl_0_6 br_0_6 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c6
*+ bl_0_6 br_0_6 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c6
*+ bl_0_6 br_0_6 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c6
*+ bl_0_6 br_0_6 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c6
*+ bl_0_6 br_0_6 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c6
*+ bl_0_6 br_0_6 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c6
*+ bl_0_6 br_0_6 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c6
*+ bl_0_6 br_0_6 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c6
*+ bl_0_6 br_0_6 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c6
*+ bl_0_6 br_0_6 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c6
*+ bl_0_6 br_0_6 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c6
*+ bl_0_6 br_0_6 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c6
*+ bl_0_6 br_0_6 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c6
*+ bl_0_6 br_0_6 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c6
*+ bl_0_6 br_0_6 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c6
*+ bl_0_6 br_0_6 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c6
*+ bl_0_6 br_0_6 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c6
*+ bl_0_6 br_0_6 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c6
*+ bl_0_6 br_0_6 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c6
*+ bl_0_6 br_0_6 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c6
*+ bl_0_6 br_0_6 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c6
*+ bl_0_6 br_0_6 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c6
*+ bl_0_6 br_0_6 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c6
*+ bl_0_6 br_0_6 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c6
*+ bl_0_6 br_0_6 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c6
*+ bl_0_6 br_0_6 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c6
*+ bl_0_6 br_0_6 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c6
*+ bl_0_6 br_0_6 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c6
*+ bl_0_6 br_0_6 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c6
*+ bl_0_6 br_0_6 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c6
*+ bl_0_6 br_0_6 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c6
*+ bl_0_6 br_0_6 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c6
*+ bl_0_6 br_0_6 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c6
*+ bl_0_6 br_0_6 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c6
*+ bl_0_6 br_0_6 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c6
*+ bl_0_6 br_0_6 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c6
*+ bl_0_6 br_0_6 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c6
*+ bl_0_6 br_0_6 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c6
*+ bl_0_6 br_0_6 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c6
*+ bl_0_6 br_0_6 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c6
*+ bl_0_6 br_0_6 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c6
*+ bl_0_6 br_0_6 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c6
*+ bl_0_6 br_0_6 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c6
*+ bl_0_6 br_0_6 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c6
*+ bl_0_6 br_0_6 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c6
*+ bl_0_6 br_0_6 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c6
*+ bl_0_6 br_0_6 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c6
*+ bl_0_6 br_0_6 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c6
*+ bl_0_6 br_0_6 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c6
*+ bl_0_6 br_0_6 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c6
*+ bl_0_6 br_0_6 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c6
*+ bl_0_6 br_0_6 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c6
*+ bl_0_6 br_0_6 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c6
*+ bl_0_6 br_0_6 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c6
*+ bl_0_6 br_0_6 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c6
*+ bl_0_6 br_0_6 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c6
*+ bl_0_6 br_0_6 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c6
*+ bl_0_6 br_0_6 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c6
*+ bl_0_6 br_0_6 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c6
*+ bl_0_6 br_0_6 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c6
*+ bl_0_6 br_0_6 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c6
*+ bl_0_6 br_0_6 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c6
*+ bl_0_6 br_0_6 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c6
*+ bl_0_6 br_0_6 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c6
*+ bl_0_6 br_0_6 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c6
*+ bl_0_6 br_0_6 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c6
*+ bl_0_6 br_0_6 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c6
*+ bl_0_6 br_0_6 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c6
*+ bl_0_6 br_0_6 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c6
*+ bl_0_6 br_0_6 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c6
*+ bl_0_6 br_0_6 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c6
*+ bl_0_6 br_0_6 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c6
*+ bl_0_6 br_0_6 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c6
*+ bl_0_6 br_0_6 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c6
*+ bl_0_6 br_0_6 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c6
*+ bl_0_6 br_0_6 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c6
*+ bl_0_6 br_0_6 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c6
*+ bl_0_6 br_0_6 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c6
*+ bl_0_6 br_0_6 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c6
*+ bl_0_6 br_0_6 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c6
*+ bl_0_6 br_0_6 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c6
*+ bl_0_6 br_0_6 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c6
*+ bl_0_6 br_0_6 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c6
*+ bl_0_6 br_0_6 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c6
*+ bl_0_6 br_0_6 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c6
*+ bl_0_6 br_0_6 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c6
*+ bl_0_6 br_0_6 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c6
*+ bl_0_6 br_0_6 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c6
*+ bl_0_6 br_0_6 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c6
*+ bl_0_6 br_0_6 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c6
*+ bl_0_6 br_0_6 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c6
*+ bl_0_6 br_0_6 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c6
*+ bl_0_6 br_0_6 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c6
*+ bl_0_6 br_0_6 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c6
*+ bl_0_6 br_0_6 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c6
*+ bl_0_6 br_0_6 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c6
*+ bl_0_6 br_0_6 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c6
*+ bl_0_6 br_0_6 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c6
*+ bl_0_6 br_0_6 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c6
*+ bl_0_6 br_0_6 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c6
*+ bl_0_6 br_0_6 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c6
*+ bl_0_6 br_0_6 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c6
*+ bl_0_6 br_0_6 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c6
*+ bl_0_6 br_0_6 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c6
*+ bl_0_6 br_0_6 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c6
*+ bl_0_6 br_0_6 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c6
*+ bl_0_6 br_0_6 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c6
*+ bl_0_6 br_0_6 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c6
*+ bl_0_6 br_0_6 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c6
*+ bl_0_6 br_0_6 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c6
*+ bl_0_6 br_0_6 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c6
*+ bl_0_6 br_0_6 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c6
*+ bl_0_6 br_0_6 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c6
*+ bl_0_6 br_0_6 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c6
+ bl_0_6 br_0_6 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c7
+ bl_0_7 br_0_7 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c7
*+ bl_0_7 br_0_7 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c7
*+ bl_0_7 br_0_7 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c7
*+ bl_0_7 br_0_7 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c7
*+ bl_0_7 br_0_7 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c7
*+ bl_0_7 br_0_7 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c7
*+ bl_0_7 br_0_7 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c7
*+ bl_0_7 br_0_7 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c7
*+ bl_0_7 br_0_7 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c7
*+ bl_0_7 br_0_7 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c7
*+ bl_0_7 br_0_7 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c7
*+ bl_0_7 br_0_7 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c7
*+ bl_0_7 br_0_7 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c7
*+ bl_0_7 br_0_7 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c7
*+ bl_0_7 br_0_7 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c7
*+ bl_0_7 br_0_7 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c7
*+ bl_0_7 br_0_7 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c7
*+ bl_0_7 br_0_7 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c7
*+ bl_0_7 br_0_7 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c7
*+ bl_0_7 br_0_7 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c7
*+ bl_0_7 br_0_7 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c7
*+ bl_0_7 br_0_7 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c7
*+ bl_0_7 br_0_7 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c7
*+ bl_0_7 br_0_7 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c7
*+ bl_0_7 br_0_7 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c7
*+ bl_0_7 br_0_7 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c7
*+ bl_0_7 br_0_7 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c7
*+ bl_0_7 br_0_7 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c7
*+ bl_0_7 br_0_7 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c7
*+ bl_0_7 br_0_7 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c7
*+ bl_0_7 br_0_7 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c7
*+ bl_0_7 br_0_7 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c7
*+ bl_0_7 br_0_7 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c7
*+ bl_0_7 br_0_7 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c7
*+ bl_0_7 br_0_7 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c7
*+ bl_0_7 br_0_7 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c7
*+ bl_0_7 br_0_7 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c7
*+ bl_0_7 br_0_7 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c7
*+ bl_0_7 br_0_7 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c7
*+ bl_0_7 br_0_7 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c7
*+ bl_0_7 br_0_7 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c7
*+ bl_0_7 br_0_7 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c7
*+ bl_0_7 br_0_7 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c7
*+ bl_0_7 br_0_7 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c7
*+ bl_0_7 br_0_7 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c7
*+ bl_0_7 br_0_7 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c7
*+ bl_0_7 br_0_7 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c7
*+ bl_0_7 br_0_7 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c7
*+ bl_0_7 br_0_7 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c7
*+ bl_0_7 br_0_7 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c7
*+ bl_0_7 br_0_7 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c7
*+ bl_0_7 br_0_7 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c7
*+ bl_0_7 br_0_7 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c7
*+ bl_0_7 br_0_7 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c7
*+ bl_0_7 br_0_7 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c7
*+ bl_0_7 br_0_7 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c7
*+ bl_0_7 br_0_7 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c7
*+ bl_0_7 br_0_7 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c7
*+ bl_0_7 br_0_7 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c7
*+ bl_0_7 br_0_7 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c7
*+ bl_0_7 br_0_7 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c7
*+ bl_0_7 br_0_7 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c7
*+ bl_0_7 br_0_7 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c7
*+ bl_0_7 br_0_7 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c7
*+ bl_0_7 br_0_7 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c7
*+ bl_0_7 br_0_7 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c7
*+ bl_0_7 br_0_7 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c7
*+ bl_0_7 br_0_7 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c7
*+ bl_0_7 br_0_7 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c7
*+ bl_0_7 br_0_7 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c7
*+ bl_0_7 br_0_7 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c7
*+ bl_0_7 br_0_7 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c7
*+ bl_0_7 br_0_7 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c7
*+ bl_0_7 br_0_7 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c7
*+ bl_0_7 br_0_7 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c7
*+ bl_0_7 br_0_7 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c7
*+ bl_0_7 br_0_7 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c7
*+ bl_0_7 br_0_7 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c7
*+ bl_0_7 br_0_7 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c7
*+ bl_0_7 br_0_7 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c7
*+ bl_0_7 br_0_7 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c7
*+ bl_0_7 br_0_7 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c7
*+ bl_0_7 br_0_7 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c7
*+ bl_0_7 br_0_7 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c7
*+ bl_0_7 br_0_7 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c7
*+ bl_0_7 br_0_7 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c7
*+ bl_0_7 br_0_7 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c7
*+ bl_0_7 br_0_7 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c7
*+ bl_0_7 br_0_7 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c7
*+ bl_0_7 br_0_7 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c7
*+ bl_0_7 br_0_7 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c7
*+ bl_0_7 br_0_7 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c7
*+ bl_0_7 br_0_7 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c7
*+ bl_0_7 br_0_7 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c7
*+ bl_0_7 br_0_7 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c7
*+ bl_0_7 br_0_7 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c7
*+ bl_0_7 br_0_7 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c7
*+ bl_0_7 br_0_7 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c7
*+ bl_0_7 br_0_7 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c7
*+ bl_0_7 br_0_7 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c7
*+ bl_0_7 br_0_7 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c7
*+ bl_0_7 br_0_7 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c7
*+ bl_0_7 br_0_7 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c7
*+ bl_0_7 br_0_7 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c7
*+ bl_0_7 br_0_7 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c7
*+ bl_0_7 br_0_7 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c7
*+ bl_0_7 br_0_7 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c7
*+ bl_0_7 br_0_7 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c7
*+ bl_0_7 br_0_7 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c7
*+ bl_0_7 br_0_7 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c7
*+ bl_0_7 br_0_7 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c7
*+ bl_0_7 br_0_7 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c7
*+ bl_0_7 br_0_7 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c7
*+ bl_0_7 br_0_7 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c7
*+ bl_0_7 br_0_7 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c7
*+ bl_0_7 br_0_7 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c7
*+ bl_0_7 br_0_7 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c7
*+ bl_0_7 br_0_7 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c7
*+ bl_0_7 br_0_7 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c7
*+ bl_0_7 br_0_7 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c7
*+ bl_0_7 br_0_7 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c7
*+ bl_0_7 br_0_7 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c7
*+ bl_0_7 br_0_7 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c7
*+ bl_0_7 br_0_7 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c7
*+ bl_0_7 br_0_7 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c7
*+ bl_0_7 br_0_7 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c7
*+ bl_0_7 br_0_7 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c7
+ bl_0_7 br_0_7 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c8
+ bl_0_8 br_0_8 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c8
*+ bl_0_8 br_0_8 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c8
*+ bl_0_8 br_0_8 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c8
*+ bl_0_8 br_0_8 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c8
*+ bl_0_8 br_0_8 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c8
*+ bl_0_8 br_0_8 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c8
*+ bl_0_8 br_0_8 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c8
*+ bl_0_8 br_0_8 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c8
*+ bl_0_8 br_0_8 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c8
*+ bl_0_8 br_0_8 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c8
*+ bl_0_8 br_0_8 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c8
*+ bl_0_8 br_0_8 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c8
*+ bl_0_8 br_0_8 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c8
*+ bl_0_8 br_0_8 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c8
*+ bl_0_8 br_0_8 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c8
*+ bl_0_8 br_0_8 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c8
*+ bl_0_8 br_0_8 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c8
*+ bl_0_8 br_0_8 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c8
*+ bl_0_8 br_0_8 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c8
*+ bl_0_8 br_0_8 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c8
*+ bl_0_8 br_0_8 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c8
*+ bl_0_8 br_0_8 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c8
*+ bl_0_8 br_0_8 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c8
*+ bl_0_8 br_0_8 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c8
*+ bl_0_8 br_0_8 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c8
*+ bl_0_8 br_0_8 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c8
*+ bl_0_8 br_0_8 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c8
*+ bl_0_8 br_0_8 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c8
*+ bl_0_8 br_0_8 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c8
*+ bl_0_8 br_0_8 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c8
*+ bl_0_8 br_0_8 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c8
*+ bl_0_8 br_0_8 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c8
*+ bl_0_8 br_0_8 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c8
*+ bl_0_8 br_0_8 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c8
*+ bl_0_8 br_0_8 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c8
*+ bl_0_8 br_0_8 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c8
*+ bl_0_8 br_0_8 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c8
*+ bl_0_8 br_0_8 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c8
*+ bl_0_8 br_0_8 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c8
*+ bl_0_8 br_0_8 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c8
*+ bl_0_8 br_0_8 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c8
*+ bl_0_8 br_0_8 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c8
*+ bl_0_8 br_0_8 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c8
*+ bl_0_8 br_0_8 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c8
*+ bl_0_8 br_0_8 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c8
*+ bl_0_8 br_0_8 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c8
*+ bl_0_8 br_0_8 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c8
*+ bl_0_8 br_0_8 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c8
*+ bl_0_8 br_0_8 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c8
*+ bl_0_8 br_0_8 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c8
*+ bl_0_8 br_0_8 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c8
*+ bl_0_8 br_0_8 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c8
*+ bl_0_8 br_0_8 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c8
*+ bl_0_8 br_0_8 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c8
*+ bl_0_8 br_0_8 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c8
*+ bl_0_8 br_0_8 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c8
*+ bl_0_8 br_0_8 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c8
*+ bl_0_8 br_0_8 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c8
*+ bl_0_8 br_0_8 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c8
*+ bl_0_8 br_0_8 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c8
*+ bl_0_8 br_0_8 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c8
*+ bl_0_8 br_0_8 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c8
*+ bl_0_8 br_0_8 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c8
*+ bl_0_8 br_0_8 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c8
*+ bl_0_8 br_0_8 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c8
*+ bl_0_8 br_0_8 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c8
*+ bl_0_8 br_0_8 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c8
*+ bl_0_8 br_0_8 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c8
*+ bl_0_8 br_0_8 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c8
*+ bl_0_8 br_0_8 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c8
*+ bl_0_8 br_0_8 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c8
*+ bl_0_8 br_0_8 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c8
*+ bl_0_8 br_0_8 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c8
*+ bl_0_8 br_0_8 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c8
*+ bl_0_8 br_0_8 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c8
*+ bl_0_8 br_0_8 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c8
*+ bl_0_8 br_0_8 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c8
*+ bl_0_8 br_0_8 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c8
*+ bl_0_8 br_0_8 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c8
*+ bl_0_8 br_0_8 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c8
*+ bl_0_8 br_0_8 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c8
*+ bl_0_8 br_0_8 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c8
*+ bl_0_8 br_0_8 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c8
*+ bl_0_8 br_0_8 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c8
*+ bl_0_8 br_0_8 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c8
*+ bl_0_8 br_0_8 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c8
*+ bl_0_8 br_0_8 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c8
*+ bl_0_8 br_0_8 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c8
*+ bl_0_8 br_0_8 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c8
*+ bl_0_8 br_0_8 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c8
*+ bl_0_8 br_0_8 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c8
*+ bl_0_8 br_0_8 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c8
*+ bl_0_8 br_0_8 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c8
*+ bl_0_8 br_0_8 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c8
*+ bl_0_8 br_0_8 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c8
*+ bl_0_8 br_0_8 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c8
*+ bl_0_8 br_0_8 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c8
*+ bl_0_8 br_0_8 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c8
*+ bl_0_8 br_0_8 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c8
*+ bl_0_8 br_0_8 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c8
*+ bl_0_8 br_0_8 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c8
*+ bl_0_8 br_0_8 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c8
*+ bl_0_8 br_0_8 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c8
*+ bl_0_8 br_0_8 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c8
*+ bl_0_8 br_0_8 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c8
*+ bl_0_8 br_0_8 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c8
*+ bl_0_8 br_0_8 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c8
*+ bl_0_8 br_0_8 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c8
*+ bl_0_8 br_0_8 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c8
*+ bl_0_8 br_0_8 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c8
*+ bl_0_8 br_0_8 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c8
*+ bl_0_8 br_0_8 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c8
*+ bl_0_8 br_0_8 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c8
*+ bl_0_8 br_0_8 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c8
*+ bl_0_8 br_0_8 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c8
*+ bl_0_8 br_0_8 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c8
*+ bl_0_8 br_0_8 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c8
*+ bl_0_8 br_0_8 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c8
*+ bl_0_8 br_0_8 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c8
*+ bl_0_8 br_0_8 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c8
*+ bl_0_8 br_0_8 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c8
*+ bl_0_8 br_0_8 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c8
*+ bl_0_8 br_0_8 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c8
*+ bl_0_8 br_0_8 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c8
*+ bl_0_8 br_0_8 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c8
*+ bl_0_8 br_0_8 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c8
*+ bl_0_8 br_0_8 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c8
+ bl_0_8 br_0_8 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c9
+ bl_0_9 br_0_9 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c9
*+ bl_0_9 br_0_9 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c9
*+ bl_0_9 br_0_9 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c9
*+ bl_0_9 br_0_9 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c9
*+ bl_0_9 br_0_9 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c9
*+ bl_0_9 br_0_9 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c9
*+ bl_0_9 br_0_9 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c9
*+ bl_0_9 br_0_9 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c9
*+ bl_0_9 br_0_9 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c9
*+ bl_0_9 br_0_9 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c9
*+ bl_0_9 br_0_9 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c9
*+ bl_0_9 br_0_9 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c9
*+ bl_0_9 br_0_9 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c9
*+ bl_0_9 br_0_9 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c9
*+ bl_0_9 br_0_9 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c9
*+ bl_0_9 br_0_9 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c9
*+ bl_0_9 br_0_9 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c9
*+ bl_0_9 br_0_9 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c9
*+ bl_0_9 br_0_9 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c9
*+ bl_0_9 br_0_9 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c9
*+ bl_0_9 br_0_9 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c9
*+ bl_0_9 br_0_9 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c9
*+ bl_0_9 br_0_9 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c9
*+ bl_0_9 br_0_9 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c9
*+ bl_0_9 br_0_9 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c9
*+ bl_0_9 br_0_9 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c9
*+ bl_0_9 br_0_9 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c9
*+ bl_0_9 br_0_9 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c9
*+ bl_0_9 br_0_9 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c9
*+ bl_0_9 br_0_9 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c9
*+ bl_0_9 br_0_9 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c9
*+ bl_0_9 br_0_9 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c9
*+ bl_0_9 br_0_9 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c9
*+ bl_0_9 br_0_9 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c9
*+ bl_0_9 br_0_9 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c9
*+ bl_0_9 br_0_9 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c9
*+ bl_0_9 br_0_9 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c9
*+ bl_0_9 br_0_9 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c9
*+ bl_0_9 br_0_9 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c9
*+ bl_0_9 br_0_9 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c9
*+ bl_0_9 br_0_9 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c9
*+ bl_0_9 br_0_9 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c9
*+ bl_0_9 br_0_9 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c9
*+ bl_0_9 br_0_9 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c9
*+ bl_0_9 br_0_9 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c9
*+ bl_0_9 br_0_9 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c9
*+ bl_0_9 br_0_9 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c9
*+ bl_0_9 br_0_9 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c9
*+ bl_0_9 br_0_9 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c9
*+ bl_0_9 br_0_9 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c9
*+ bl_0_9 br_0_9 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c9
*+ bl_0_9 br_0_9 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c9
*+ bl_0_9 br_0_9 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c9
*+ bl_0_9 br_0_9 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c9
*+ bl_0_9 br_0_9 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c9
*+ bl_0_9 br_0_9 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c9
*+ bl_0_9 br_0_9 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c9
*+ bl_0_9 br_0_9 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c9
*+ bl_0_9 br_0_9 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c9
*+ bl_0_9 br_0_9 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c9
*+ bl_0_9 br_0_9 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c9
*+ bl_0_9 br_0_9 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c9
*+ bl_0_9 br_0_9 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c9
*+ bl_0_9 br_0_9 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c9
*+ bl_0_9 br_0_9 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c9
*+ bl_0_9 br_0_9 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c9
*+ bl_0_9 br_0_9 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c9
*+ bl_0_9 br_0_9 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c9
*+ bl_0_9 br_0_9 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c9
*+ bl_0_9 br_0_9 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c9
*+ bl_0_9 br_0_9 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c9
*+ bl_0_9 br_0_9 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c9
*+ bl_0_9 br_0_9 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c9
*+ bl_0_9 br_0_9 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c9
*+ bl_0_9 br_0_9 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c9
*+ bl_0_9 br_0_9 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c9
*+ bl_0_9 br_0_9 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c9
*+ bl_0_9 br_0_9 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c9
*+ bl_0_9 br_0_9 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c9
*+ bl_0_9 br_0_9 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c9
*+ bl_0_9 br_0_9 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c9
*+ bl_0_9 br_0_9 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c9
*+ bl_0_9 br_0_9 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c9
*+ bl_0_9 br_0_9 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c9
*+ bl_0_9 br_0_9 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c9
*+ bl_0_9 br_0_9 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c9
*+ bl_0_9 br_0_9 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c9
*+ bl_0_9 br_0_9 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c9
*+ bl_0_9 br_0_9 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c9
*+ bl_0_9 br_0_9 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c9
*+ bl_0_9 br_0_9 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c9
*+ bl_0_9 br_0_9 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c9
*+ bl_0_9 br_0_9 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c9
*+ bl_0_9 br_0_9 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c9
*+ bl_0_9 br_0_9 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c9
*+ bl_0_9 br_0_9 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c9
*+ bl_0_9 br_0_9 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c9
*+ bl_0_9 br_0_9 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c9
*+ bl_0_9 br_0_9 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c9
*+ bl_0_9 br_0_9 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c9
*+ bl_0_9 br_0_9 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c9
*+ bl_0_9 br_0_9 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c9
*+ bl_0_9 br_0_9 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c9
*+ bl_0_9 br_0_9 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c9
*+ bl_0_9 br_0_9 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c9
*+ bl_0_9 br_0_9 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c9
*+ bl_0_9 br_0_9 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c9
*+ bl_0_9 br_0_9 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c9
*+ bl_0_9 br_0_9 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c9
*+ bl_0_9 br_0_9 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c9
*+ bl_0_9 br_0_9 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c9
*+ bl_0_9 br_0_9 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c9
*+ bl_0_9 br_0_9 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c9
*+ bl_0_9 br_0_9 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c9
*+ bl_0_9 br_0_9 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c9
*+ bl_0_9 br_0_9 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c9
*+ bl_0_9 br_0_9 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c9
*+ bl_0_9 br_0_9 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c9
*+ bl_0_9 br_0_9 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c9
*+ bl_0_9 br_0_9 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c9
*+ bl_0_9 br_0_9 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c9
*+ bl_0_9 br_0_9 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c9
*+ bl_0_9 br_0_9 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c9
*+ bl_0_9 br_0_9 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c9
*+ bl_0_9 br_0_9 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c9
*+ bl_0_9 br_0_9 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c9
*+ bl_0_9 br_0_9 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c9
+ bl_0_9 br_0_9 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c10
+ bl_0_10 br_0_10 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c10
*+ bl_0_10 br_0_10 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c10
*+ bl_0_10 br_0_10 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c10
*+ bl_0_10 br_0_10 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c10
*+ bl_0_10 br_0_10 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c10
*+ bl_0_10 br_0_10 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c10
*+ bl_0_10 br_0_10 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c10
*+ bl_0_10 br_0_10 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c10
*+ bl_0_10 br_0_10 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c10
*+ bl_0_10 br_0_10 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c10
*+ bl_0_10 br_0_10 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c10
*+ bl_0_10 br_0_10 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c10
*+ bl_0_10 br_0_10 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c10
*+ bl_0_10 br_0_10 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c10
*+ bl_0_10 br_0_10 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c10
*+ bl_0_10 br_0_10 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c10
*+ bl_0_10 br_0_10 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c10
*+ bl_0_10 br_0_10 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c10
*+ bl_0_10 br_0_10 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c10
*+ bl_0_10 br_0_10 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c10
*+ bl_0_10 br_0_10 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c10
*+ bl_0_10 br_0_10 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c10
*+ bl_0_10 br_0_10 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c10
*+ bl_0_10 br_0_10 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c10
*+ bl_0_10 br_0_10 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c10
*+ bl_0_10 br_0_10 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c10
*+ bl_0_10 br_0_10 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c10
*+ bl_0_10 br_0_10 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c10
*+ bl_0_10 br_0_10 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c10
*+ bl_0_10 br_0_10 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c10
*+ bl_0_10 br_0_10 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c10
*+ bl_0_10 br_0_10 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c10
*+ bl_0_10 br_0_10 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c10
*+ bl_0_10 br_0_10 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c10
*+ bl_0_10 br_0_10 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c10
*+ bl_0_10 br_0_10 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c10
*+ bl_0_10 br_0_10 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c10
*+ bl_0_10 br_0_10 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c10
*+ bl_0_10 br_0_10 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c10
*+ bl_0_10 br_0_10 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c10
*+ bl_0_10 br_0_10 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c10
*+ bl_0_10 br_0_10 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c10
*+ bl_0_10 br_0_10 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c10
*+ bl_0_10 br_0_10 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c10
*+ bl_0_10 br_0_10 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c10
*+ bl_0_10 br_0_10 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c10
*+ bl_0_10 br_0_10 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c10
*+ bl_0_10 br_0_10 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c10
*+ bl_0_10 br_0_10 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c10
*+ bl_0_10 br_0_10 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c10
*+ bl_0_10 br_0_10 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c10
*+ bl_0_10 br_0_10 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c10
*+ bl_0_10 br_0_10 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c10
*+ bl_0_10 br_0_10 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c10
*+ bl_0_10 br_0_10 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c10
*+ bl_0_10 br_0_10 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c10
*+ bl_0_10 br_0_10 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c10
*+ bl_0_10 br_0_10 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c10
*+ bl_0_10 br_0_10 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c10
*+ bl_0_10 br_0_10 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c10
*+ bl_0_10 br_0_10 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c10
*+ bl_0_10 br_0_10 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c10
*+ bl_0_10 br_0_10 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c10
*+ bl_0_10 br_0_10 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c10
*+ bl_0_10 br_0_10 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c10
*+ bl_0_10 br_0_10 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c10
*+ bl_0_10 br_0_10 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c10
*+ bl_0_10 br_0_10 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c10
*+ bl_0_10 br_0_10 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c10
*+ bl_0_10 br_0_10 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c10
*+ bl_0_10 br_0_10 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c10
*+ bl_0_10 br_0_10 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c10
*+ bl_0_10 br_0_10 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c10
*+ bl_0_10 br_0_10 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c10
*+ bl_0_10 br_0_10 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c10
*+ bl_0_10 br_0_10 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c10
*+ bl_0_10 br_0_10 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c10
*+ bl_0_10 br_0_10 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c10
*+ bl_0_10 br_0_10 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c10
*+ bl_0_10 br_0_10 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c10
*+ bl_0_10 br_0_10 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c10
*+ bl_0_10 br_0_10 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c10
*+ bl_0_10 br_0_10 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c10
*+ bl_0_10 br_0_10 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c10
*+ bl_0_10 br_0_10 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c10
*+ bl_0_10 br_0_10 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c10
*+ bl_0_10 br_0_10 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c10
*+ bl_0_10 br_0_10 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c10
*+ bl_0_10 br_0_10 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c10
*+ bl_0_10 br_0_10 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c10
*+ bl_0_10 br_0_10 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c10
*+ bl_0_10 br_0_10 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c10
*+ bl_0_10 br_0_10 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c10
*+ bl_0_10 br_0_10 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c10
*+ bl_0_10 br_0_10 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c10
*+ bl_0_10 br_0_10 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c10
*+ bl_0_10 br_0_10 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c10
*+ bl_0_10 br_0_10 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c10
*+ bl_0_10 br_0_10 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c10
*+ bl_0_10 br_0_10 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c10
*+ bl_0_10 br_0_10 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c10
*+ bl_0_10 br_0_10 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c10
*+ bl_0_10 br_0_10 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c10
*+ bl_0_10 br_0_10 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c10
*+ bl_0_10 br_0_10 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c10
*+ bl_0_10 br_0_10 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c10
*+ bl_0_10 br_0_10 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c10
*+ bl_0_10 br_0_10 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c10
*+ bl_0_10 br_0_10 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c10
*+ bl_0_10 br_0_10 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c10
*+ bl_0_10 br_0_10 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c10
*+ bl_0_10 br_0_10 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c10
*+ bl_0_10 br_0_10 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c10
*+ bl_0_10 br_0_10 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c10
*+ bl_0_10 br_0_10 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c10
*+ bl_0_10 br_0_10 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c10
*+ bl_0_10 br_0_10 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c10
*+ bl_0_10 br_0_10 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c10
*+ bl_0_10 br_0_10 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c10
*+ bl_0_10 br_0_10 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c10
*+ bl_0_10 br_0_10 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c10
*+ bl_0_10 br_0_10 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c10
*+ bl_0_10 br_0_10 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c10
*+ bl_0_10 br_0_10 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c10
*+ bl_0_10 br_0_10 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c10
*+ bl_0_10 br_0_10 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c10
*+ bl_0_10 br_0_10 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c10
+ bl_0_10 br_0_10 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c11
+ bl_0_11 br_0_11 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c11
*+ bl_0_11 br_0_11 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c11
*+ bl_0_11 br_0_11 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c11
*+ bl_0_11 br_0_11 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c11
*+ bl_0_11 br_0_11 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c11
*+ bl_0_11 br_0_11 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c11
*+ bl_0_11 br_0_11 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c11
*+ bl_0_11 br_0_11 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c11
*+ bl_0_11 br_0_11 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c11
*+ bl_0_11 br_0_11 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c11
*+ bl_0_11 br_0_11 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c11
*+ bl_0_11 br_0_11 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c11
*+ bl_0_11 br_0_11 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c11
*+ bl_0_11 br_0_11 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c11
*+ bl_0_11 br_0_11 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c11
*+ bl_0_11 br_0_11 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c11
*+ bl_0_11 br_0_11 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c11
*+ bl_0_11 br_0_11 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c11
*+ bl_0_11 br_0_11 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c11
*+ bl_0_11 br_0_11 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c11
*+ bl_0_11 br_0_11 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c11
*+ bl_0_11 br_0_11 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c11
*+ bl_0_11 br_0_11 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c11
*+ bl_0_11 br_0_11 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c11
*+ bl_0_11 br_0_11 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c11
*+ bl_0_11 br_0_11 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c11
*+ bl_0_11 br_0_11 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c11
*+ bl_0_11 br_0_11 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c11
*+ bl_0_11 br_0_11 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c11
*+ bl_0_11 br_0_11 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c11
*+ bl_0_11 br_0_11 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c11
*+ bl_0_11 br_0_11 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c11
*+ bl_0_11 br_0_11 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c11
*+ bl_0_11 br_0_11 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c11
*+ bl_0_11 br_0_11 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c11
*+ bl_0_11 br_0_11 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c11
*+ bl_0_11 br_0_11 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c11
*+ bl_0_11 br_0_11 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c11
*+ bl_0_11 br_0_11 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c11
*+ bl_0_11 br_0_11 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c11
*+ bl_0_11 br_0_11 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c11
*+ bl_0_11 br_0_11 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c11
*+ bl_0_11 br_0_11 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c11
*+ bl_0_11 br_0_11 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c11
*+ bl_0_11 br_0_11 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c11
*+ bl_0_11 br_0_11 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c11
*+ bl_0_11 br_0_11 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c11
*+ bl_0_11 br_0_11 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c11
*+ bl_0_11 br_0_11 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c11
*+ bl_0_11 br_0_11 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c11
*+ bl_0_11 br_0_11 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c11
*+ bl_0_11 br_0_11 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c11
*+ bl_0_11 br_0_11 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c11
*+ bl_0_11 br_0_11 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c11
*+ bl_0_11 br_0_11 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c11
*+ bl_0_11 br_0_11 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c11
*+ bl_0_11 br_0_11 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c11
*+ bl_0_11 br_0_11 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c11
*+ bl_0_11 br_0_11 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c11
*+ bl_0_11 br_0_11 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c11
*+ bl_0_11 br_0_11 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c11
*+ bl_0_11 br_0_11 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c11
*+ bl_0_11 br_0_11 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c11
*+ bl_0_11 br_0_11 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c11
*+ bl_0_11 br_0_11 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c11
*+ bl_0_11 br_0_11 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c11
*+ bl_0_11 br_0_11 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c11
*+ bl_0_11 br_0_11 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c11
*+ bl_0_11 br_0_11 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c11
*+ bl_0_11 br_0_11 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c11
*+ bl_0_11 br_0_11 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c11
*+ bl_0_11 br_0_11 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c11
*+ bl_0_11 br_0_11 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c11
*+ bl_0_11 br_0_11 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c11
*+ bl_0_11 br_0_11 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c11
*+ bl_0_11 br_0_11 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c11
*+ bl_0_11 br_0_11 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c11
*+ bl_0_11 br_0_11 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c11
*+ bl_0_11 br_0_11 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c11
*+ bl_0_11 br_0_11 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c11
*+ bl_0_11 br_0_11 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c11
*+ bl_0_11 br_0_11 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c11
*+ bl_0_11 br_0_11 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c11
*+ bl_0_11 br_0_11 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c11
*+ bl_0_11 br_0_11 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c11
*+ bl_0_11 br_0_11 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c11
*+ bl_0_11 br_0_11 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c11
*+ bl_0_11 br_0_11 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c11
*+ bl_0_11 br_0_11 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c11
*+ bl_0_11 br_0_11 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c11
*+ bl_0_11 br_0_11 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c11
*+ bl_0_11 br_0_11 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c11
*+ bl_0_11 br_0_11 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c11
*+ bl_0_11 br_0_11 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c11
*+ bl_0_11 br_0_11 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c11
*+ bl_0_11 br_0_11 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c11
*+ bl_0_11 br_0_11 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c11
*+ bl_0_11 br_0_11 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c11
*+ bl_0_11 br_0_11 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c11
*+ bl_0_11 br_0_11 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c11
*+ bl_0_11 br_0_11 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c11
*+ bl_0_11 br_0_11 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c11
*+ bl_0_11 br_0_11 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c11
*+ bl_0_11 br_0_11 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c11
*+ bl_0_11 br_0_11 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c11
*+ bl_0_11 br_0_11 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c11
*+ bl_0_11 br_0_11 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c11
*+ bl_0_11 br_0_11 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c11
*+ bl_0_11 br_0_11 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c11
*+ bl_0_11 br_0_11 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c11
*+ bl_0_11 br_0_11 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c11
*+ bl_0_11 br_0_11 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c11
*+ bl_0_11 br_0_11 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c11
*+ bl_0_11 br_0_11 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c11
*+ bl_0_11 br_0_11 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c11
*+ bl_0_11 br_0_11 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c11
*+ bl_0_11 br_0_11 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c11
*+ bl_0_11 br_0_11 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c11
*+ bl_0_11 br_0_11 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c11
*+ bl_0_11 br_0_11 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c11
*+ bl_0_11 br_0_11 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c11
*+ bl_0_11 br_0_11 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c11
*+ bl_0_11 br_0_11 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c11
*+ bl_0_11 br_0_11 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c11
*+ bl_0_11 br_0_11 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c11
*+ bl_0_11 br_0_11 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c11
*+ bl_0_11 br_0_11 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c11
+ bl_0_11 br_0_11 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c12
+ bl_0_12 br_0_12 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c12
*+ bl_0_12 br_0_12 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c12
*+ bl_0_12 br_0_12 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c12
*+ bl_0_12 br_0_12 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c12
*+ bl_0_12 br_0_12 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c12
*+ bl_0_12 br_0_12 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c12
*+ bl_0_12 br_0_12 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c12
*+ bl_0_12 br_0_12 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c12
*+ bl_0_12 br_0_12 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c12
*+ bl_0_12 br_0_12 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c12
*+ bl_0_12 br_0_12 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c12
*+ bl_0_12 br_0_12 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c12
*+ bl_0_12 br_0_12 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c12
*+ bl_0_12 br_0_12 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c12
*+ bl_0_12 br_0_12 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c12
*+ bl_0_12 br_0_12 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c12
*+ bl_0_12 br_0_12 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c12
*+ bl_0_12 br_0_12 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c12
*+ bl_0_12 br_0_12 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c12
*+ bl_0_12 br_0_12 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c12
*+ bl_0_12 br_0_12 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c12
*+ bl_0_12 br_0_12 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c12
*+ bl_0_12 br_0_12 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c12
*+ bl_0_12 br_0_12 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c12
*+ bl_0_12 br_0_12 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c12
*+ bl_0_12 br_0_12 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c12
*+ bl_0_12 br_0_12 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c12
*+ bl_0_12 br_0_12 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c12
*+ bl_0_12 br_0_12 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c12
*+ bl_0_12 br_0_12 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c12
*+ bl_0_12 br_0_12 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c12
*+ bl_0_12 br_0_12 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c12
*+ bl_0_12 br_0_12 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c12
*+ bl_0_12 br_0_12 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c12
*+ bl_0_12 br_0_12 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c12
*+ bl_0_12 br_0_12 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c12
*+ bl_0_12 br_0_12 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c12
*+ bl_0_12 br_0_12 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c12
*+ bl_0_12 br_0_12 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c12
*+ bl_0_12 br_0_12 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c12
*+ bl_0_12 br_0_12 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c12
*+ bl_0_12 br_0_12 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c12
*+ bl_0_12 br_0_12 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c12
*+ bl_0_12 br_0_12 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c12
*+ bl_0_12 br_0_12 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c12
*+ bl_0_12 br_0_12 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c12
*+ bl_0_12 br_0_12 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c12
*+ bl_0_12 br_0_12 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c12
*+ bl_0_12 br_0_12 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c12
*+ bl_0_12 br_0_12 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c12
*+ bl_0_12 br_0_12 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c12
*+ bl_0_12 br_0_12 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c12
*+ bl_0_12 br_0_12 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c12
*+ bl_0_12 br_0_12 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c12
*+ bl_0_12 br_0_12 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c12
*+ bl_0_12 br_0_12 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c12
*+ bl_0_12 br_0_12 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c12
*+ bl_0_12 br_0_12 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c12
*+ bl_0_12 br_0_12 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c12
*+ bl_0_12 br_0_12 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c12
*+ bl_0_12 br_0_12 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c12
*+ bl_0_12 br_0_12 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c12
*+ bl_0_12 br_0_12 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c12
*+ bl_0_12 br_0_12 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c12
*+ bl_0_12 br_0_12 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c12
*+ bl_0_12 br_0_12 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c12
*+ bl_0_12 br_0_12 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c12
*+ bl_0_12 br_0_12 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c12
*+ bl_0_12 br_0_12 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c12
*+ bl_0_12 br_0_12 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c12
*+ bl_0_12 br_0_12 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c12
*+ bl_0_12 br_0_12 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c12
*+ bl_0_12 br_0_12 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c12
*+ bl_0_12 br_0_12 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c12
*+ bl_0_12 br_0_12 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c12
*+ bl_0_12 br_0_12 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c12
*+ bl_0_12 br_0_12 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c12
*+ bl_0_12 br_0_12 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c12
*+ bl_0_12 br_0_12 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c12
*+ bl_0_12 br_0_12 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c12
*+ bl_0_12 br_0_12 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c12
*+ bl_0_12 br_0_12 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c12
*+ bl_0_12 br_0_12 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c12
*+ bl_0_12 br_0_12 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c12
*+ bl_0_12 br_0_12 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c12
*+ bl_0_12 br_0_12 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c12
*+ bl_0_12 br_0_12 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c12
*+ bl_0_12 br_0_12 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c12
*+ bl_0_12 br_0_12 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c12
*+ bl_0_12 br_0_12 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c12
*+ bl_0_12 br_0_12 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c12
*+ bl_0_12 br_0_12 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c12
*+ bl_0_12 br_0_12 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c12
*+ bl_0_12 br_0_12 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c12
*+ bl_0_12 br_0_12 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c12
*+ bl_0_12 br_0_12 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c12
*+ bl_0_12 br_0_12 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c12
*+ bl_0_12 br_0_12 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c12
*+ bl_0_12 br_0_12 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c12
*+ bl_0_12 br_0_12 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c12
*+ bl_0_12 br_0_12 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c12
*+ bl_0_12 br_0_12 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c12
*+ bl_0_12 br_0_12 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c12
*+ bl_0_12 br_0_12 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c12
*+ bl_0_12 br_0_12 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c12
*+ bl_0_12 br_0_12 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c12
*+ bl_0_12 br_0_12 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c12
*+ bl_0_12 br_0_12 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c12
*+ bl_0_12 br_0_12 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c12
*+ bl_0_12 br_0_12 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c12
*+ bl_0_12 br_0_12 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c12
*+ bl_0_12 br_0_12 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c12
*+ bl_0_12 br_0_12 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c12
*+ bl_0_12 br_0_12 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c12
*+ bl_0_12 br_0_12 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c12
*+ bl_0_12 br_0_12 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c12
*+ bl_0_12 br_0_12 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c12
*+ bl_0_12 br_0_12 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c12
*+ bl_0_12 br_0_12 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c12
*+ bl_0_12 br_0_12 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c12
*+ bl_0_12 br_0_12 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c12
*+ bl_0_12 br_0_12 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c12
*+ bl_0_12 br_0_12 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c12
*+ bl_0_12 br_0_12 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c12
*+ bl_0_12 br_0_12 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c12
*+ bl_0_12 br_0_12 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c12
*+ bl_0_12 br_0_12 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c12
+ bl_0_12 br_0_12 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c13
+ bl_0_13 br_0_13 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c13
*+ bl_0_13 br_0_13 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c13
*+ bl_0_13 br_0_13 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c13
*+ bl_0_13 br_0_13 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c13
*+ bl_0_13 br_0_13 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c13
*+ bl_0_13 br_0_13 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c13
*+ bl_0_13 br_0_13 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c13
*+ bl_0_13 br_0_13 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c13
*+ bl_0_13 br_0_13 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c13
*+ bl_0_13 br_0_13 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c13
*+ bl_0_13 br_0_13 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c13
*+ bl_0_13 br_0_13 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c13
*+ bl_0_13 br_0_13 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c13
*+ bl_0_13 br_0_13 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c13
*+ bl_0_13 br_0_13 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c13
*+ bl_0_13 br_0_13 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c13
*+ bl_0_13 br_0_13 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c13
*+ bl_0_13 br_0_13 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c13
*+ bl_0_13 br_0_13 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c13
*+ bl_0_13 br_0_13 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c13
*+ bl_0_13 br_0_13 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c13
*+ bl_0_13 br_0_13 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c13
*+ bl_0_13 br_0_13 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c13
*+ bl_0_13 br_0_13 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c13
*+ bl_0_13 br_0_13 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c13
*+ bl_0_13 br_0_13 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c13
*+ bl_0_13 br_0_13 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c13
*+ bl_0_13 br_0_13 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c13
*+ bl_0_13 br_0_13 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c13
*+ bl_0_13 br_0_13 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c13
*+ bl_0_13 br_0_13 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c13
*+ bl_0_13 br_0_13 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c13
*+ bl_0_13 br_0_13 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c13
*+ bl_0_13 br_0_13 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c13
*+ bl_0_13 br_0_13 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c13
*+ bl_0_13 br_0_13 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c13
*+ bl_0_13 br_0_13 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c13
*+ bl_0_13 br_0_13 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c13
*+ bl_0_13 br_0_13 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c13
*+ bl_0_13 br_0_13 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c13
*+ bl_0_13 br_0_13 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c13
*+ bl_0_13 br_0_13 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c13
*+ bl_0_13 br_0_13 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c13
*+ bl_0_13 br_0_13 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c13
*+ bl_0_13 br_0_13 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c13
*+ bl_0_13 br_0_13 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c13
*+ bl_0_13 br_0_13 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c13
*+ bl_0_13 br_0_13 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c13
*+ bl_0_13 br_0_13 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c13
*+ bl_0_13 br_0_13 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c13
*+ bl_0_13 br_0_13 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c13
*+ bl_0_13 br_0_13 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c13
*+ bl_0_13 br_0_13 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c13
*+ bl_0_13 br_0_13 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c13
*+ bl_0_13 br_0_13 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c13
*+ bl_0_13 br_0_13 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c13
*+ bl_0_13 br_0_13 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c13
*+ bl_0_13 br_0_13 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c13
*+ bl_0_13 br_0_13 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c13
*+ bl_0_13 br_0_13 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c13
*+ bl_0_13 br_0_13 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c13
*+ bl_0_13 br_0_13 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c13
*+ bl_0_13 br_0_13 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c13
*+ bl_0_13 br_0_13 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c13
*+ bl_0_13 br_0_13 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c13
*+ bl_0_13 br_0_13 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c13
*+ bl_0_13 br_0_13 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c13
*+ bl_0_13 br_0_13 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c13
*+ bl_0_13 br_0_13 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c13
*+ bl_0_13 br_0_13 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c13
*+ bl_0_13 br_0_13 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c13
*+ bl_0_13 br_0_13 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c13
*+ bl_0_13 br_0_13 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c13
*+ bl_0_13 br_0_13 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c13
*+ bl_0_13 br_0_13 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c13
*+ bl_0_13 br_0_13 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c13
*+ bl_0_13 br_0_13 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c13
*+ bl_0_13 br_0_13 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c13
*+ bl_0_13 br_0_13 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c13
*+ bl_0_13 br_0_13 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c13
*+ bl_0_13 br_0_13 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c13
*+ bl_0_13 br_0_13 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c13
*+ bl_0_13 br_0_13 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c13
*+ bl_0_13 br_0_13 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c13
*+ bl_0_13 br_0_13 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c13
*+ bl_0_13 br_0_13 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c13
*+ bl_0_13 br_0_13 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c13
*+ bl_0_13 br_0_13 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c13
*+ bl_0_13 br_0_13 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c13
*+ bl_0_13 br_0_13 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c13
*+ bl_0_13 br_0_13 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c13
*+ bl_0_13 br_0_13 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c13
*+ bl_0_13 br_0_13 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c13
*+ bl_0_13 br_0_13 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c13
*+ bl_0_13 br_0_13 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c13
*+ bl_0_13 br_0_13 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c13
*+ bl_0_13 br_0_13 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c13
*+ bl_0_13 br_0_13 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c13
*+ bl_0_13 br_0_13 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c13
*+ bl_0_13 br_0_13 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c13
*+ bl_0_13 br_0_13 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c13
*+ bl_0_13 br_0_13 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c13
*+ bl_0_13 br_0_13 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c13
*+ bl_0_13 br_0_13 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c13
*+ bl_0_13 br_0_13 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c13
*+ bl_0_13 br_0_13 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c13
*+ bl_0_13 br_0_13 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c13
*+ bl_0_13 br_0_13 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c13
*+ bl_0_13 br_0_13 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c13
*+ bl_0_13 br_0_13 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c13
*+ bl_0_13 br_0_13 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c13
*+ bl_0_13 br_0_13 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c13
*+ bl_0_13 br_0_13 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c13
*+ bl_0_13 br_0_13 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c13
*+ bl_0_13 br_0_13 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c13
*+ bl_0_13 br_0_13 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c13
*+ bl_0_13 br_0_13 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c13
*+ bl_0_13 br_0_13 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c13
*+ bl_0_13 br_0_13 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c13
*+ bl_0_13 br_0_13 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c13
*+ bl_0_13 br_0_13 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c13
*+ bl_0_13 br_0_13 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c13
*+ bl_0_13 br_0_13 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c13
*+ bl_0_13 br_0_13 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c13
*+ bl_0_13 br_0_13 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c13
*+ bl_0_13 br_0_13 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c13
*+ bl_0_13 br_0_13 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c13
+ bl_0_13 br_0_13 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c14
+ bl_0_14 br_0_14 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c14
*+ bl_0_14 br_0_14 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c14
*+ bl_0_14 br_0_14 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c14
*+ bl_0_14 br_0_14 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c14
*+ bl_0_14 br_0_14 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c14
*+ bl_0_14 br_0_14 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c14
*+ bl_0_14 br_0_14 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c14
*+ bl_0_14 br_0_14 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c14
*+ bl_0_14 br_0_14 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c14
*+ bl_0_14 br_0_14 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c14
*+ bl_0_14 br_0_14 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c14
*+ bl_0_14 br_0_14 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c14
*+ bl_0_14 br_0_14 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c14
*+ bl_0_14 br_0_14 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c14
*+ bl_0_14 br_0_14 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c14
*+ bl_0_14 br_0_14 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c14
*+ bl_0_14 br_0_14 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c14
*+ bl_0_14 br_0_14 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c14
*+ bl_0_14 br_0_14 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c14
*+ bl_0_14 br_0_14 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c14
*+ bl_0_14 br_0_14 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c14
*+ bl_0_14 br_0_14 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c14
*+ bl_0_14 br_0_14 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c14
*+ bl_0_14 br_0_14 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c14
*+ bl_0_14 br_0_14 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c14
*+ bl_0_14 br_0_14 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c14
*+ bl_0_14 br_0_14 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c14
*+ bl_0_14 br_0_14 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c14
*+ bl_0_14 br_0_14 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c14
*+ bl_0_14 br_0_14 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c14
*+ bl_0_14 br_0_14 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c14
*+ bl_0_14 br_0_14 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c14
*+ bl_0_14 br_0_14 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c14
*+ bl_0_14 br_0_14 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c14
*+ bl_0_14 br_0_14 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c14
*+ bl_0_14 br_0_14 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c14
*+ bl_0_14 br_0_14 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c14
*+ bl_0_14 br_0_14 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c14
*+ bl_0_14 br_0_14 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c14
*+ bl_0_14 br_0_14 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c14
*+ bl_0_14 br_0_14 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c14
*+ bl_0_14 br_0_14 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c14
*+ bl_0_14 br_0_14 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c14
*+ bl_0_14 br_0_14 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c14
*+ bl_0_14 br_0_14 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c14
*+ bl_0_14 br_0_14 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c14
*+ bl_0_14 br_0_14 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c14
*+ bl_0_14 br_0_14 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c14
*+ bl_0_14 br_0_14 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c14
*+ bl_0_14 br_0_14 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c14
*+ bl_0_14 br_0_14 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c14
*+ bl_0_14 br_0_14 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c14
*+ bl_0_14 br_0_14 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c14
*+ bl_0_14 br_0_14 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c14
*+ bl_0_14 br_0_14 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c14
*+ bl_0_14 br_0_14 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c14
*+ bl_0_14 br_0_14 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c14
*+ bl_0_14 br_0_14 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c14
*+ bl_0_14 br_0_14 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c14
*+ bl_0_14 br_0_14 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c14
*+ bl_0_14 br_0_14 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c14
*+ bl_0_14 br_0_14 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c14
*+ bl_0_14 br_0_14 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c14
*+ bl_0_14 br_0_14 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c14
*+ bl_0_14 br_0_14 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c14
*+ bl_0_14 br_0_14 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c14
*+ bl_0_14 br_0_14 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c14
*+ bl_0_14 br_0_14 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c14
*+ bl_0_14 br_0_14 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c14
*+ bl_0_14 br_0_14 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c14
*+ bl_0_14 br_0_14 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c14
*+ bl_0_14 br_0_14 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c14
*+ bl_0_14 br_0_14 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c14
*+ bl_0_14 br_0_14 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c14
*+ bl_0_14 br_0_14 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c14
*+ bl_0_14 br_0_14 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c14
*+ bl_0_14 br_0_14 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c14
*+ bl_0_14 br_0_14 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c14
*+ bl_0_14 br_0_14 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c14
*+ bl_0_14 br_0_14 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c14
*+ bl_0_14 br_0_14 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c14
*+ bl_0_14 br_0_14 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c14
*+ bl_0_14 br_0_14 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c14
*+ bl_0_14 br_0_14 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c14
*+ bl_0_14 br_0_14 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c14
*+ bl_0_14 br_0_14 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c14
*+ bl_0_14 br_0_14 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c14
*+ bl_0_14 br_0_14 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c14
*+ bl_0_14 br_0_14 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c14
*+ bl_0_14 br_0_14 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c14
*+ bl_0_14 br_0_14 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c14
*+ bl_0_14 br_0_14 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c14
*+ bl_0_14 br_0_14 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c14
*+ bl_0_14 br_0_14 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c14
*+ bl_0_14 br_0_14 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c14
*+ bl_0_14 br_0_14 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c14
*+ bl_0_14 br_0_14 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c14
*+ bl_0_14 br_0_14 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c14
*+ bl_0_14 br_0_14 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c14
*+ bl_0_14 br_0_14 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c14
*+ bl_0_14 br_0_14 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c14
*+ bl_0_14 br_0_14 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c14
*+ bl_0_14 br_0_14 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c14
*+ bl_0_14 br_0_14 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c14
*+ bl_0_14 br_0_14 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c14
*+ bl_0_14 br_0_14 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c14
*+ bl_0_14 br_0_14 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c14
*+ bl_0_14 br_0_14 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c14
*+ bl_0_14 br_0_14 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c14
*+ bl_0_14 br_0_14 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c14
*+ bl_0_14 br_0_14 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c14
*+ bl_0_14 br_0_14 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c14
*+ bl_0_14 br_0_14 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c14
*+ bl_0_14 br_0_14 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c14
*+ bl_0_14 br_0_14 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c14
*+ bl_0_14 br_0_14 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c14
*+ bl_0_14 br_0_14 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c14
*+ bl_0_14 br_0_14 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c14
*+ bl_0_14 br_0_14 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c14
*+ bl_0_14 br_0_14 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c14
*+ bl_0_14 br_0_14 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c14
*+ bl_0_14 br_0_14 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c14
*+ bl_0_14 br_0_14 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c14
*+ bl_0_14 br_0_14 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c14
*+ bl_0_14 br_0_14 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c14
*+ bl_0_14 br_0_14 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c14
*+ bl_0_14 br_0_14 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c14
+ bl_0_14 br_0_14 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c15
+ bl_0_15 br_0_15 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c15
*+ bl_0_15 br_0_15 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c15
*+ bl_0_15 br_0_15 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c15
*+ bl_0_15 br_0_15 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c15
*+ bl_0_15 br_0_15 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c15
*+ bl_0_15 br_0_15 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c15
*+ bl_0_15 br_0_15 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c15
*+ bl_0_15 br_0_15 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c15
*+ bl_0_15 br_0_15 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c15
*+ bl_0_15 br_0_15 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c15
*+ bl_0_15 br_0_15 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c15
*+ bl_0_15 br_0_15 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c15
*+ bl_0_15 br_0_15 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c15
*+ bl_0_15 br_0_15 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c15
*+ bl_0_15 br_0_15 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c15
*+ bl_0_15 br_0_15 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c15
*+ bl_0_15 br_0_15 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c15
*+ bl_0_15 br_0_15 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c15
*+ bl_0_15 br_0_15 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c15
*+ bl_0_15 br_0_15 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c15
*+ bl_0_15 br_0_15 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c15
*+ bl_0_15 br_0_15 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c15
*+ bl_0_15 br_0_15 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c15
*+ bl_0_15 br_0_15 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c15
*+ bl_0_15 br_0_15 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c15
*+ bl_0_15 br_0_15 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c15
*+ bl_0_15 br_0_15 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c15
*+ bl_0_15 br_0_15 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c15
*+ bl_0_15 br_0_15 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c15
*+ bl_0_15 br_0_15 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c15
*+ bl_0_15 br_0_15 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c15
*+ bl_0_15 br_0_15 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c15
*+ bl_0_15 br_0_15 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c15
*+ bl_0_15 br_0_15 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c15
*+ bl_0_15 br_0_15 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c15
*+ bl_0_15 br_0_15 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c15
*+ bl_0_15 br_0_15 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c15
*+ bl_0_15 br_0_15 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c15
*+ bl_0_15 br_0_15 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c15
*+ bl_0_15 br_0_15 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c15
*+ bl_0_15 br_0_15 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c15
*+ bl_0_15 br_0_15 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c15
*+ bl_0_15 br_0_15 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c15
*+ bl_0_15 br_0_15 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c15
*+ bl_0_15 br_0_15 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c15
*+ bl_0_15 br_0_15 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c15
*+ bl_0_15 br_0_15 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c15
*+ bl_0_15 br_0_15 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c15
*+ bl_0_15 br_0_15 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c15
*+ bl_0_15 br_0_15 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c15
*+ bl_0_15 br_0_15 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c15
*+ bl_0_15 br_0_15 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c15
*+ bl_0_15 br_0_15 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c15
*+ bl_0_15 br_0_15 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c15
*+ bl_0_15 br_0_15 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c15
*+ bl_0_15 br_0_15 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c15
*+ bl_0_15 br_0_15 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c15
*+ bl_0_15 br_0_15 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c15
*+ bl_0_15 br_0_15 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c15
*+ bl_0_15 br_0_15 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c15
*+ bl_0_15 br_0_15 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c15
*+ bl_0_15 br_0_15 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c15
*+ bl_0_15 br_0_15 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c15
*+ bl_0_15 br_0_15 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c15
*+ bl_0_15 br_0_15 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c15
*+ bl_0_15 br_0_15 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c15
*+ bl_0_15 br_0_15 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c15
*+ bl_0_15 br_0_15 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c15
*+ bl_0_15 br_0_15 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c15
*+ bl_0_15 br_0_15 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c15
*+ bl_0_15 br_0_15 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c15
*+ bl_0_15 br_0_15 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c15
*+ bl_0_15 br_0_15 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c15
*+ bl_0_15 br_0_15 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c15
*+ bl_0_15 br_0_15 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c15
*+ bl_0_15 br_0_15 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c15
*+ bl_0_15 br_0_15 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c15
*+ bl_0_15 br_0_15 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c15
*+ bl_0_15 br_0_15 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c15
*+ bl_0_15 br_0_15 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c15
*+ bl_0_15 br_0_15 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c15
*+ bl_0_15 br_0_15 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c15
*+ bl_0_15 br_0_15 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c15
*+ bl_0_15 br_0_15 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c15
*+ bl_0_15 br_0_15 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c15
*+ bl_0_15 br_0_15 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c15
*+ bl_0_15 br_0_15 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c15
*+ bl_0_15 br_0_15 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c15
*+ bl_0_15 br_0_15 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c15
*+ bl_0_15 br_0_15 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c15
*+ bl_0_15 br_0_15 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c15
*+ bl_0_15 br_0_15 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c15
*+ bl_0_15 br_0_15 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c15
*+ bl_0_15 br_0_15 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c15
*+ bl_0_15 br_0_15 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c15
*+ bl_0_15 br_0_15 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c15
*+ bl_0_15 br_0_15 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c15
*+ bl_0_15 br_0_15 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c15
*+ bl_0_15 br_0_15 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c15
*+ bl_0_15 br_0_15 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c15
*+ bl_0_15 br_0_15 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c15
*+ bl_0_15 br_0_15 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c15
*+ bl_0_15 br_0_15 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c15
*+ bl_0_15 br_0_15 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c15
*+ bl_0_15 br_0_15 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c15
*+ bl_0_15 br_0_15 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c15
*+ bl_0_15 br_0_15 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c15
*+ bl_0_15 br_0_15 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c15
*+ bl_0_15 br_0_15 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c15
*+ bl_0_15 br_0_15 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c15
*+ bl_0_15 br_0_15 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c15
*+ bl_0_15 br_0_15 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c15
*+ bl_0_15 br_0_15 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c15
*+ bl_0_15 br_0_15 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c15
*+ bl_0_15 br_0_15 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c15
*+ bl_0_15 br_0_15 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c15
*+ bl_0_15 br_0_15 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c15
*+ bl_0_15 br_0_15 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c15
*+ bl_0_15 br_0_15 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c15
*+ bl_0_15 br_0_15 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c15
*+ bl_0_15 br_0_15 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c15
*+ bl_0_15 br_0_15 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c15
*+ bl_0_15 br_0_15 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c15
*+ bl_0_15 br_0_15 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c15
*+ bl_0_15 br_0_15 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c15
*+ bl_0_15 br_0_15 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c15
*+ bl_0_15 br_0_15 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c15
+ bl_0_15 br_0_15 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c16
+ bl_0_16 br_0_16 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c16
*+ bl_0_16 br_0_16 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c16
*+ bl_0_16 br_0_16 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c16
*+ bl_0_16 br_0_16 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c16
*+ bl_0_16 br_0_16 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c16
*+ bl_0_16 br_0_16 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c16
*+ bl_0_16 br_0_16 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c16
*+ bl_0_16 br_0_16 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c16
*+ bl_0_16 br_0_16 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c16
*+ bl_0_16 br_0_16 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c16
*+ bl_0_16 br_0_16 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c16
*+ bl_0_16 br_0_16 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c16
*+ bl_0_16 br_0_16 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c16
*+ bl_0_16 br_0_16 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c16
*+ bl_0_16 br_0_16 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c16
*+ bl_0_16 br_0_16 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c16
*+ bl_0_16 br_0_16 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c16
*+ bl_0_16 br_0_16 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c16
*+ bl_0_16 br_0_16 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c16
*+ bl_0_16 br_0_16 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c16
*+ bl_0_16 br_0_16 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c16
*+ bl_0_16 br_0_16 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c16
*+ bl_0_16 br_0_16 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c16
*+ bl_0_16 br_0_16 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c16
*+ bl_0_16 br_0_16 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c16
*+ bl_0_16 br_0_16 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c16
*+ bl_0_16 br_0_16 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c16
*+ bl_0_16 br_0_16 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c16
*+ bl_0_16 br_0_16 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c16
*+ bl_0_16 br_0_16 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c16
*+ bl_0_16 br_0_16 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c16
*+ bl_0_16 br_0_16 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c16
*+ bl_0_16 br_0_16 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c16
*+ bl_0_16 br_0_16 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c16
*+ bl_0_16 br_0_16 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c16
*+ bl_0_16 br_0_16 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c16
*+ bl_0_16 br_0_16 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c16
*+ bl_0_16 br_0_16 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c16
*+ bl_0_16 br_0_16 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c16
*+ bl_0_16 br_0_16 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c16
*+ bl_0_16 br_0_16 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c16
*+ bl_0_16 br_0_16 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c16
*+ bl_0_16 br_0_16 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c16
*+ bl_0_16 br_0_16 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c16
*+ bl_0_16 br_0_16 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c16
*+ bl_0_16 br_0_16 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c16
*+ bl_0_16 br_0_16 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c16
*+ bl_0_16 br_0_16 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c16
*+ bl_0_16 br_0_16 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c16
*+ bl_0_16 br_0_16 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c16
*+ bl_0_16 br_0_16 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c16
*+ bl_0_16 br_0_16 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c16
*+ bl_0_16 br_0_16 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c16
*+ bl_0_16 br_0_16 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c16
*+ bl_0_16 br_0_16 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c16
*+ bl_0_16 br_0_16 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c16
*+ bl_0_16 br_0_16 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c16
*+ bl_0_16 br_0_16 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c16
*+ bl_0_16 br_0_16 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c16
*+ bl_0_16 br_0_16 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c16
*+ bl_0_16 br_0_16 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c16
*+ bl_0_16 br_0_16 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c16
*+ bl_0_16 br_0_16 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c16
*+ bl_0_16 br_0_16 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c16
*+ bl_0_16 br_0_16 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c16
*+ bl_0_16 br_0_16 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c16
*+ bl_0_16 br_0_16 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c16
*+ bl_0_16 br_0_16 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c16
*+ bl_0_16 br_0_16 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c16
*+ bl_0_16 br_0_16 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c16
*+ bl_0_16 br_0_16 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c16
*+ bl_0_16 br_0_16 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c16
*+ bl_0_16 br_0_16 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c16
*+ bl_0_16 br_0_16 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c16
*+ bl_0_16 br_0_16 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c16
*+ bl_0_16 br_0_16 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c16
*+ bl_0_16 br_0_16 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c16
*+ bl_0_16 br_0_16 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c16
*+ bl_0_16 br_0_16 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c16
*+ bl_0_16 br_0_16 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c16
*+ bl_0_16 br_0_16 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c16
*+ bl_0_16 br_0_16 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c16
*+ bl_0_16 br_0_16 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c16
*+ bl_0_16 br_0_16 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c16
*+ bl_0_16 br_0_16 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c16
*+ bl_0_16 br_0_16 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c16
*+ bl_0_16 br_0_16 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c16
*+ bl_0_16 br_0_16 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c16
*+ bl_0_16 br_0_16 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c16
*+ bl_0_16 br_0_16 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c16
*+ bl_0_16 br_0_16 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c16
*+ bl_0_16 br_0_16 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c16
*+ bl_0_16 br_0_16 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c16
*+ bl_0_16 br_0_16 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c16
*+ bl_0_16 br_0_16 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c16
*+ bl_0_16 br_0_16 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c16
*+ bl_0_16 br_0_16 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c16
*+ bl_0_16 br_0_16 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c16
*+ bl_0_16 br_0_16 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c16
*+ bl_0_16 br_0_16 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c16
*+ bl_0_16 br_0_16 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c16
*+ bl_0_16 br_0_16 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c16
*+ bl_0_16 br_0_16 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c16
*+ bl_0_16 br_0_16 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c16
*+ bl_0_16 br_0_16 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c16
*+ bl_0_16 br_0_16 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c16
*+ bl_0_16 br_0_16 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c16
*+ bl_0_16 br_0_16 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c16
*+ bl_0_16 br_0_16 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c16
*+ bl_0_16 br_0_16 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c16
*+ bl_0_16 br_0_16 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c16
*+ bl_0_16 br_0_16 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c16
*+ bl_0_16 br_0_16 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c16
*+ bl_0_16 br_0_16 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c16
*+ bl_0_16 br_0_16 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c16
*+ bl_0_16 br_0_16 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c16
*+ bl_0_16 br_0_16 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c16
*+ bl_0_16 br_0_16 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c16
*+ bl_0_16 br_0_16 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c16
*+ bl_0_16 br_0_16 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c16
*+ bl_0_16 br_0_16 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c16
*+ bl_0_16 br_0_16 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c16
*+ bl_0_16 br_0_16 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c16
*+ bl_0_16 br_0_16 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c16
*+ bl_0_16 br_0_16 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c16
*+ bl_0_16 br_0_16 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c16
*+ bl_0_16 br_0_16 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c16
+ bl_0_16 br_0_16 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c17
+ bl_0_17 br_0_17 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c17
*+ bl_0_17 br_0_17 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c17
*+ bl_0_17 br_0_17 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c17
*+ bl_0_17 br_0_17 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c17
*+ bl_0_17 br_0_17 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c17
*+ bl_0_17 br_0_17 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c17
*+ bl_0_17 br_0_17 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c17
*+ bl_0_17 br_0_17 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c17
*+ bl_0_17 br_0_17 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c17
*+ bl_0_17 br_0_17 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c17
*+ bl_0_17 br_0_17 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c17
*+ bl_0_17 br_0_17 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c17
*+ bl_0_17 br_0_17 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c17
*+ bl_0_17 br_0_17 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c17
*+ bl_0_17 br_0_17 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c17
*+ bl_0_17 br_0_17 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c17
*+ bl_0_17 br_0_17 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c17
*+ bl_0_17 br_0_17 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c17
*+ bl_0_17 br_0_17 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c17
*+ bl_0_17 br_0_17 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c17
*+ bl_0_17 br_0_17 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c17
*+ bl_0_17 br_0_17 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c17
*+ bl_0_17 br_0_17 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c17
*+ bl_0_17 br_0_17 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c17
*+ bl_0_17 br_0_17 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c17
*+ bl_0_17 br_0_17 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c17
*+ bl_0_17 br_0_17 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c17
*+ bl_0_17 br_0_17 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c17
*+ bl_0_17 br_0_17 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c17
*+ bl_0_17 br_0_17 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c17
*+ bl_0_17 br_0_17 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c17
*+ bl_0_17 br_0_17 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c17
*+ bl_0_17 br_0_17 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c17
*+ bl_0_17 br_0_17 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c17
*+ bl_0_17 br_0_17 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c17
*+ bl_0_17 br_0_17 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c17
*+ bl_0_17 br_0_17 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c17
*+ bl_0_17 br_0_17 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c17
*+ bl_0_17 br_0_17 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c17
*+ bl_0_17 br_0_17 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c17
*+ bl_0_17 br_0_17 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c17
*+ bl_0_17 br_0_17 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c17
*+ bl_0_17 br_0_17 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c17
*+ bl_0_17 br_0_17 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c17
*+ bl_0_17 br_0_17 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c17
*+ bl_0_17 br_0_17 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c17
*+ bl_0_17 br_0_17 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c17
*+ bl_0_17 br_0_17 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c17
*+ bl_0_17 br_0_17 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c17
*+ bl_0_17 br_0_17 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c17
*+ bl_0_17 br_0_17 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c17
*+ bl_0_17 br_0_17 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c17
*+ bl_0_17 br_0_17 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c17
*+ bl_0_17 br_0_17 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c17
*+ bl_0_17 br_0_17 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c17
*+ bl_0_17 br_0_17 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c17
*+ bl_0_17 br_0_17 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c17
*+ bl_0_17 br_0_17 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c17
*+ bl_0_17 br_0_17 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c17
*+ bl_0_17 br_0_17 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c17
*+ bl_0_17 br_0_17 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c17
*+ bl_0_17 br_0_17 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c17
*+ bl_0_17 br_0_17 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c17
*+ bl_0_17 br_0_17 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c17
*+ bl_0_17 br_0_17 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c17
*+ bl_0_17 br_0_17 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c17
*+ bl_0_17 br_0_17 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c17
*+ bl_0_17 br_0_17 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c17
*+ bl_0_17 br_0_17 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c17
*+ bl_0_17 br_0_17 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c17
*+ bl_0_17 br_0_17 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c17
*+ bl_0_17 br_0_17 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c17
*+ bl_0_17 br_0_17 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c17
*+ bl_0_17 br_0_17 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c17
*+ bl_0_17 br_0_17 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c17
*+ bl_0_17 br_0_17 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c17
*+ bl_0_17 br_0_17 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c17
*+ bl_0_17 br_0_17 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c17
*+ bl_0_17 br_0_17 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c17
*+ bl_0_17 br_0_17 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c17
*+ bl_0_17 br_0_17 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c17
*+ bl_0_17 br_0_17 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c17
*+ bl_0_17 br_0_17 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c17
*+ bl_0_17 br_0_17 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c17
*+ bl_0_17 br_0_17 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c17
*+ bl_0_17 br_0_17 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c17
*+ bl_0_17 br_0_17 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c17
*+ bl_0_17 br_0_17 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c17
*+ bl_0_17 br_0_17 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c17
*+ bl_0_17 br_0_17 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c17
*+ bl_0_17 br_0_17 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c17
*+ bl_0_17 br_0_17 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c17
*+ bl_0_17 br_0_17 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c17
*+ bl_0_17 br_0_17 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c17
*+ bl_0_17 br_0_17 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c17
*+ bl_0_17 br_0_17 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c17
*+ bl_0_17 br_0_17 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c17
*+ bl_0_17 br_0_17 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c17
*+ bl_0_17 br_0_17 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c17
*+ bl_0_17 br_0_17 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c17
*+ bl_0_17 br_0_17 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c17
*+ bl_0_17 br_0_17 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c17
*+ bl_0_17 br_0_17 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c17
*+ bl_0_17 br_0_17 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c17
*+ bl_0_17 br_0_17 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c17
*+ bl_0_17 br_0_17 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c17
*+ bl_0_17 br_0_17 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c17
*+ bl_0_17 br_0_17 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c17
*+ bl_0_17 br_0_17 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c17
*+ bl_0_17 br_0_17 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c17
*+ bl_0_17 br_0_17 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c17
*+ bl_0_17 br_0_17 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c17
*+ bl_0_17 br_0_17 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c17
*+ bl_0_17 br_0_17 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c17
*+ bl_0_17 br_0_17 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c17
*+ bl_0_17 br_0_17 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c17
*+ bl_0_17 br_0_17 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c17
*+ bl_0_17 br_0_17 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c17
*+ bl_0_17 br_0_17 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c17
*+ bl_0_17 br_0_17 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c17
*+ bl_0_17 br_0_17 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c17
*+ bl_0_17 br_0_17 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c17
*+ bl_0_17 br_0_17 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c17
*+ bl_0_17 br_0_17 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c17
*+ bl_0_17 br_0_17 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c17
*+ bl_0_17 br_0_17 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c17
*+ bl_0_17 br_0_17 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c17
+ bl_0_17 br_0_17 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c18
+ bl_0_18 br_0_18 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c18
*+ bl_0_18 br_0_18 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c18
*+ bl_0_18 br_0_18 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c18
*+ bl_0_18 br_0_18 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c18
*+ bl_0_18 br_0_18 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c18
*+ bl_0_18 br_0_18 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c18
*+ bl_0_18 br_0_18 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c18
*+ bl_0_18 br_0_18 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c18
*+ bl_0_18 br_0_18 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c18
*+ bl_0_18 br_0_18 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c18
*+ bl_0_18 br_0_18 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c18
*+ bl_0_18 br_0_18 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c18
*+ bl_0_18 br_0_18 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c18
*+ bl_0_18 br_0_18 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c18
*+ bl_0_18 br_0_18 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c18
*+ bl_0_18 br_0_18 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c18
*+ bl_0_18 br_0_18 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c18
*+ bl_0_18 br_0_18 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c18
*+ bl_0_18 br_0_18 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c18
*+ bl_0_18 br_0_18 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c18
*+ bl_0_18 br_0_18 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c18
*+ bl_0_18 br_0_18 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c18
*+ bl_0_18 br_0_18 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c18
*+ bl_0_18 br_0_18 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c18
*+ bl_0_18 br_0_18 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c18
*+ bl_0_18 br_0_18 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c18
*+ bl_0_18 br_0_18 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c18
*+ bl_0_18 br_0_18 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c18
*+ bl_0_18 br_0_18 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c18
*+ bl_0_18 br_0_18 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c18
*+ bl_0_18 br_0_18 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c18
*+ bl_0_18 br_0_18 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c18
*+ bl_0_18 br_0_18 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c18
*+ bl_0_18 br_0_18 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c18
*+ bl_0_18 br_0_18 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c18
*+ bl_0_18 br_0_18 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c18
*+ bl_0_18 br_0_18 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c18
*+ bl_0_18 br_0_18 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c18
*+ bl_0_18 br_0_18 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c18
*+ bl_0_18 br_0_18 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c18
*+ bl_0_18 br_0_18 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c18
*+ bl_0_18 br_0_18 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c18
*+ bl_0_18 br_0_18 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c18
*+ bl_0_18 br_0_18 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c18
*+ bl_0_18 br_0_18 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c18
*+ bl_0_18 br_0_18 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c18
*+ bl_0_18 br_0_18 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c18
*+ bl_0_18 br_0_18 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c18
*+ bl_0_18 br_0_18 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c18
*+ bl_0_18 br_0_18 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c18
*+ bl_0_18 br_0_18 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c18
*+ bl_0_18 br_0_18 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c18
*+ bl_0_18 br_0_18 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c18
*+ bl_0_18 br_0_18 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c18
*+ bl_0_18 br_0_18 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c18
*+ bl_0_18 br_0_18 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c18
*+ bl_0_18 br_0_18 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c18
*+ bl_0_18 br_0_18 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c18
*+ bl_0_18 br_0_18 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c18
*+ bl_0_18 br_0_18 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c18
*+ bl_0_18 br_0_18 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c18
*+ bl_0_18 br_0_18 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c18
*+ bl_0_18 br_0_18 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c18
*+ bl_0_18 br_0_18 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c18
*+ bl_0_18 br_0_18 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c18
*+ bl_0_18 br_0_18 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c18
*+ bl_0_18 br_0_18 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c18
*+ bl_0_18 br_0_18 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c18
*+ bl_0_18 br_0_18 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c18
*+ bl_0_18 br_0_18 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c18
*+ bl_0_18 br_0_18 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c18
*+ bl_0_18 br_0_18 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c18
*+ bl_0_18 br_0_18 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c18
*+ bl_0_18 br_0_18 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c18
*+ bl_0_18 br_0_18 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c18
*+ bl_0_18 br_0_18 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c18
*+ bl_0_18 br_0_18 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c18
*+ bl_0_18 br_0_18 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c18
*+ bl_0_18 br_0_18 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c18
*+ bl_0_18 br_0_18 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c18
*+ bl_0_18 br_0_18 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c18
*+ bl_0_18 br_0_18 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c18
*+ bl_0_18 br_0_18 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c18
*+ bl_0_18 br_0_18 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c18
*+ bl_0_18 br_0_18 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c18
*+ bl_0_18 br_0_18 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c18
*+ bl_0_18 br_0_18 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c18
*+ bl_0_18 br_0_18 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c18
*+ bl_0_18 br_0_18 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c18
*+ bl_0_18 br_0_18 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c18
*+ bl_0_18 br_0_18 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c18
*+ bl_0_18 br_0_18 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c18
*+ bl_0_18 br_0_18 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c18
*+ bl_0_18 br_0_18 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c18
*+ bl_0_18 br_0_18 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c18
*+ bl_0_18 br_0_18 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c18
*+ bl_0_18 br_0_18 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c18
*+ bl_0_18 br_0_18 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c18
*+ bl_0_18 br_0_18 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c18
*+ bl_0_18 br_0_18 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c18
*+ bl_0_18 br_0_18 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c18
*+ bl_0_18 br_0_18 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c18
*+ bl_0_18 br_0_18 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c18
*+ bl_0_18 br_0_18 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c18
*+ bl_0_18 br_0_18 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c18
*+ bl_0_18 br_0_18 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c18
*+ bl_0_18 br_0_18 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c18
*+ bl_0_18 br_0_18 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c18
*+ bl_0_18 br_0_18 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c18
*+ bl_0_18 br_0_18 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c18
*+ bl_0_18 br_0_18 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c18
*+ bl_0_18 br_0_18 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c18
*+ bl_0_18 br_0_18 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c18
*+ bl_0_18 br_0_18 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c18
*+ bl_0_18 br_0_18 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c18
*+ bl_0_18 br_0_18 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c18
*+ bl_0_18 br_0_18 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c18
*+ bl_0_18 br_0_18 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c18
*+ bl_0_18 br_0_18 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c18
*+ bl_0_18 br_0_18 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c18
*+ bl_0_18 br_0_18 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c18
*+ bl_0_18 br_0_18 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c18
*+ bl_0_18 br_0_18 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c18
*+ bl_0_18 br_0_18 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c18
*+ bl_0_18 br_0_18 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c18
*+ bl_0_18 br_0_18 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c18
*+ bl_0_18 br_0_18 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c18
+ bl_0_18 br_0_18 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c19
+ bl_0_19 br_0_19 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c19
*+ bl_0_19 br_0_19 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c19
*+ bl_0_19 br_0_19 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c19
*+ bl_0_19 br_0_19 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c19
*+ bl_0_19 br_0_19 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c19
*+ bl_0_19 br_0_19 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c19
*+ bl_0_19 br_0_19 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c19
*+ bl_0_19 br_0_19 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c19
*+ bl_0_19 br_0_19 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c19
*+ bl_0_19 br_0_19 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c19
*+ bl_0_19 br_0_19 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c19
*+ bl_0_19 br_0_19 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c19
*+ bl_0_19 br_0_19 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c19
*+ bl_0_19 br_0_19 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c19
*+ bl_0_19 br_0_19 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c19
*+ bl_0_19 br_0_19 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c19
*+ bl_0_19 br_0_19 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c19
*+ bl_0_19 br_0_19 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c19
*+ bl_0_19 br_0_19 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c19
*+ bl_0_19 br_0_19 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c19
*+ bl_0_19 br_0_19 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c19
*+ bl_0_19 br_0_19 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c19
*+ bl_0_19 br_0_19 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c19
*+ bl_0_19 br_0_19 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c19
*+ bl_0_19 br_0_19 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c19
*+ bl_0_19 br_0_19 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c19
*+ bl_0_19 br_0_19 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c19
*+ bl_0_19 br_0_19 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c19
*+ bl_0_19 br_0_19 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c19
*+ bl_0_19 br_0_19 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c19
*+ bl_0_19 br_0_19 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c19
*+ bl_0_19 br_0_19 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c19
*+ bl_0_19 br_0_19 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c19
*+ bl_0_19 br_0_19 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c19
*+ bl_0_19 br_0_19 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c19
*+ bl_0_19 br_0_19 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c19
*+ bl_0_19 br_0_19 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c19
*+ bl_0_19 br_0_19 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c19
*+ bl_0_19 br_0_19 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c19
*+ bl_0_19 br_0_19 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c19
*+ bl_0_19 br_0_19 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c19
*+ bl_0_19 br_0_19 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c19
*+ bl_0_19 br_0_19 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c19
*+ bl_0_19 br_0_19 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c19
*+ bl_0_19 br_0_19 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c19
*+ bl_0_19 br_0_19 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c19
*+ bl_0_19 br_0_19 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c19
*+ bl_0_19 br_0_19 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c19
*+ bl_0_19 br_0_19 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c19
*+ bl_0_19 br_0_19 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c19
*+ bl_0_19 br_0_19 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c19
*+ bl_0_19 br_0_19 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c19
*+ bl_0_19 br_0_19 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c19
*+ bl_0_19 br_0_19 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c19
*+ bl_0_19 br_0_19 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c19
*+ bl_0_19 br_0_19 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c19
*+ bl_0_19 br_0_19 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c19
*+ bl_0_19 br_0_19 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c19
*+ bl_0_19 br_0_19 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c19
*+ bl_0_19 br_0_19 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c19
*+ bl_0_19 br_0_19 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c19
*+ bl_0_19 br_0_19 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c19
*+ bl_0_19 br_0_19 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c19
*+ bl_0_19 br_0_19 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c19
*+ bl_0_19 br_0_19 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c19
*+ bl_0_19 br_0_19 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c19
*+ bl_0_19 br_0_19 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c19
*+ bl_0_19 br_0_19 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c19
*+ bl_0_19 br_0_19 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c19
*+ bl_0_19 br_0_19 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c19
*+ bl_0_19 br_0_19 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c19
*+ bl_0_19 br_0_19 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c19
*+ bl_0_19 br_0_19 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c19
*+ bl_0_19 br_0_19 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c19
*+ bl_0_19 br_0_19 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c19
*+ bl_0_19 br_0_19 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c19
*+ bl_0_19 br_0_19 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c19
*+ bl_0_19 br_0_19 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c19
*+ bl_0_19 br_0_19 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c19
*+ bl_0_19 br_0_19 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c19
*+ bl_0_19 br_0_19 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c19
*+ bl_0_19 br_0_19 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c19
*+ bl_0_19 br_0_19 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c19
*+ bl_0_19 br_0_19 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c19
*+ bl_0_19 br_0_19 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c19
*+ bl_0_19 br_0_19 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c19
*+ bl_0_19 br_0_19 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c19
*+ bl_0_19 br_0_19 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c19
*+ bl_0_19 br_0_19 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c19
*+ bl_0_19 br_0_19 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c19
*+ bl_0_19 br_0_19 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c19
*+ bl_0_19 br_0_19 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c19
*+ bl_0_19 br_0_19 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c19
*+ bl_0_19 br_0_19 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c19
*+ bl_0_19 br_0_19 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c19
*+ bl_0_19 br_0_19 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c19
*+ bl_0_19 br_0_19 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c19
*+ bl_0_19 br_0_19 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c19
*+ bl_0_19 br_0_19 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c19
*+ bl_0_19 br_0_19 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c19
*+ bl_0_19 br_0_19 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c19
*+ bl_0_19 br_0_19 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c19
*+ bl_0_19 br_0_19 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c19
*+ bl_0_19 br_0_19 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c19
*+ bl_0_19 br_0_19 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c19
*+ bl_0_19 br_0_19 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c19
*+ bl_0_19 br_0_19 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c19
*+ bl_0_19 br_0_19 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c19
*+ bl_0_19 br_0_19 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c19
*+ bl_0_19 br_0_19 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c19
*+ bl_0_19 br_0_19 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c19
*+ bl_0_19 br_0_19 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c19
*+ bl_0_19 br_0_19 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c19
*+ bl_0_19 br_0_19 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c19
*+ bl_0_19 br_0_19 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c19
*+ bl_0_19 br_0_19 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c19
*+ bl_0_19 br_0_19 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c19
*+ bl_0_19 br_0_19 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c19
*+ bl_0_19 br_0_19 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c19
*+ bl_0_19 br_0_19 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c19
*+ bl_0_19 br_0_19 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c19
*+ bl_0_19 br_0_19 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c19
*+ bl_0_19 br_0_19 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c19
*+ bl_0_19 br_0_19 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c19
*+ bl_0_19 br_0_19 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c19
*+ bl_0_19 br_0_19 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c19
*+ bl_0_19 br_0_19 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c19
+ bl_0_19 br_0_19 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c20
+ bl_0_20 br_0_20 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c20
*+ bl_0_20 br_0_20 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c20
*+ bl_0_20 br_0_20 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c20
*+ bl_0_20 br_0_20 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c20
*+ bl_0_20 br_0_20 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c20
*+ bl_0_20 br_0_20 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c20
*+ bl_0_20 br_0_20 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c20
*+ bl_0_20 br_0_20 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c20
*+ bl_0_20 br_0_20 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c20
*+ bl_0_20 br_0_20 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c20
*+ bl_0_20 br_0_20 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c20
*+ bl_0_20 br_0_20 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c20
*+ bl_0_20 br_0_20 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c20
*+ bl_0_20 br_0_20 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c20
*+ bl_0_20 br_0_20 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c20
*+ bl_0_20 br_0_20 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c20
*+ bl_0_20 br_0_20 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c20
*+ bl_0_20 br_0_20 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c20
*+ bl_0_20 br_0_20 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c20
*+ bl_0_20 br_0_20 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c20
*+ bl_0_20 br_0_20 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c20
*+ bl_0_20 br_0_20 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c20
*+ bl_0_20 br_0_20 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c20
*+ bl_0_20 br_0_20 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c20
*+ bl_0_20 br_0_20 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c20
*+ bl_0_20 br_0_20 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c20
*+ bl_0_20 br_0_20 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c20
*+ bl_0_20 br_0_20 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c20
*+ bl_0_20 br_0_20 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c20
*+ bl_0_20 br_0_20 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c20
*+ bl_0_20 br_0_20 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c20
*+ bl_0_20 br_0_20 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c20
*+ bl_0_20 br_0_20 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c20
*+ bl_0_20 br_0_20 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c20
*+ bl_0_20 br_0_20 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c20
*+ bl_0_20 br_0_20 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c20
*+ bl_0_20 br_0_20 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c20
*+ bl_0_20 br_0_20 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c20
*+ bl_0_20 br_0_20 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c20
*+ bl_0_20 br_0_20 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c20
*+ bl_0_20 br_0_20 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c20
*+ bl_0_20 br_0_20 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c20
*+ bl_0_20 br_0_20 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c20
*+ bl_0_20 br_0_20 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c20
*+ bl_0_20 br_0_20 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c20
*+ bl_0_20 br_0_20 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c20
*+ bl_0_20 br_0_20 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c20
*+ bl_0_20 br_0_20 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c20
*+ bl_0_20 br_0_20 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c20
*+ bl_0_20 br_0_20 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c20
*+ bl_0_20 br_0_20 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c20
*+ bl_0_20 br_0_20 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c20
*+ bl_0_20 br_0_20 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c20
*+ bl_0_20 br_0_20 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c20
*+ bl_0_20 br_0_20 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c20
*+ bl_0_20 br_0_20 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c20
*+ bl_0_20 br_0_20 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c20
*+ bl_0_20 br_0_20 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c20
*+ bl_0_20 br_0_20 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c20
*+ bl_0_20 br_0_20 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c20
*+ bl_0_20 br_0_20 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c20
*+ bl_0_20 br_0_20 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c20
*+ bl_0_20 br_0_20 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c20
*+ bl_0_20 br_0_20 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c20
*+ bl_0_20 br_0_20 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c20
*+ bl_0_20 br_0_20 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c20
*+ bl_0_20 br_0_20 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c20
*+ bl_0_20 br_0_20 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c20
*+ bl_0_20 br_0_20 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c20
*+ bl_0_20 br_0_20 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c20
*+ bl_0_20 br_0_20 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c20
*+ bl_0_20 br_0_20 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c20
*+ bl_0_20 br_0_20 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c20
*+ bl_0_20 br_0_20 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c20
*+ bl_0_20 br_0_20 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c20
*+ bl_0_20 br_0_20 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c20
*+ bl_0_20 br_0_20 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c20
*+ bl_0_20 br_0_20 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c20
*+ bl_0_20 br_0_20 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c20
*+ bl_0_20 br_0_20 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c20
*+ bl_0_20 br_0_20 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c20
*+ bl_0_20 br_0_20 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c20
*+ bl_0_20 br_0_20 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c20
*+ bl_0_20 br_0_20 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c20
*+ bl_0_20 br_0_20 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c20
*+ bl_0_20 br_0_20 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c20
*+ bl_0_20 br_0_20 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c20
*+ bl_0_20 br_0_20 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c20
*+ bl_0_20 br_0_20 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c20
*+ bl_0_20 br_0_20 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c20
*+ bl_0_20 br_0_20 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c20
*+ bl_0_20 br_0_20 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c20
*+ bl_0_20 br_0_20 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c20
*+ bl_0_20 br_0_20 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c20
*+ bl_0_20 br_0_20 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c20
*+ bl_0_20 br_0_20 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c20
*+ bl_0_20 br_0_20 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c20
*+ bl_0_20 br_0_20 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c20
*+ bl_0_20 br_0_20 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c20
*+ bl_0_20 br_0_20 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c20
*+ bl_0_20 br_0_20 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c20
*+ bl_0_20 br_0_20 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c20
*+ bl_0_20 br_0_20 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c20
*+ bl_0_20 br_0_20 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c20
*+ bl_0_20 br_0_20 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c20
*+ bl_0_20 br_0_20 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c20
*+ bl_0_20 br_0_20 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c20
*+ bl_0_20 br_0_20 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c20
*+ bl_0_20 br_0_20 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c20
*+ bl_0_20 br_0_20 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c20
*+ bl_0_20 br_0_20 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c20
*+ bl_0_20 br_0_20 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c20
*+ bl_0_20 br_0_20 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c20
*+ bl_0_20 br_0_20 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c20
*+ bl_0_20 br_0_20 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c20
*+ bl_0_20 br_0_20 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c20
*+ bl_0_20 br_0_20 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c20
*+ bl_0_20 br_0_20 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c20
*+ bl_0_20 br_0_20 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c20
*+ bl_0_20 br_0_20 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c20
*+ bl_0_20 br_0_20 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c20
*+ bl_0_20 br_0_20 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c20
*+ bl_0_20 br_0_20 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c20
*+ bl_0_20 br_0_20 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c20
*+ bl_0_20 br_0_20 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c20
*+ bl_0_20 br_0_20 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c20
*+ bl_0_20 br_0_20 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c20
+ bl_0_20 br_0_20 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c21
+ bl_0_21 br_0_21 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c21
*+ bl_0_21 br_0_21 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c21
*+ bl_0_21 br_0_21 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c21
*+ bl_0_21 br_0_21 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c21
*+ bl_0_21 br_0_21 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c21
*+ bl_0_21 br_0_21 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c21
*+ bl_0_21 br_0_21 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c21
*+ bl_0_21 br_0_21 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c21
*+ bl_0_21 br_0_21 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c21
*+ bl_0_21 br_0_21 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c21
*+ bl_0_21 br_0_21 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c21
*+ bl_0_21 br_0_21 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c21
*+ bl_0_21 br_0_21 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c21
*+ bl_0_21 br_0_21 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c21
*+ bl_0_21 br_0_21 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c21
*+ bl_0_21 br_0_21 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c21
*+ bl_0_21 br_0_21 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c21
*+ bl_0_21 br_0_21 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c21
*+ bl_0_21 br_0_21 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c21
*+ bl_0_21 br_0_21 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c21
*+ bl_0_21 br_0_21 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c21
*+ bl_0_21 br_0_21 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c21
*+ bl_0_21 br_0_21 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c21
*+ bl_0_21 br_0_21 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c21
*+ bl_0_21 br_0_21 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c21
*+ bl_0_21 br_0_21 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c21
*+ bl_0_21 br_0_21 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c21
*+ bl_0_21 br_0_21 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c21
*+ bl_0_21 br_0_21 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c21
*+ bl_0_21 br_0_21 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c21
*+ bl_0_21 br_0_21 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c21
*+ bl_0_21 br_0_21 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c21
*+ bl_0_21 br_0_21 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c21
*+ bl_0_21 br_0_21 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c21
*+ bl_0_21 br_0_21 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c21
*+ bl_0_21 br_0_21 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c21
*+ bl_0_21 br_0_21 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c21
*+ bl_0_21 br_0_21 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c21
*+ bl_0_21 br_0_21 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c21
*+ bl_0_21 br_0_21 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c21
*+ bl_0_21 br_0_21 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c21
*+ bl_0_21 br_0_21 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c21
*+ bl_0_21 br_0_21 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c21
*+ bl_0_21 br_0_21 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c21
*+ bl_0_21 br_0_21 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c21
*+ bl_0_21 br_0_21 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c21
*+ bl_0_21 br_0_21 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c21
*+ bl_0_21 br_0_21 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c21
*+ bl_0_21 br_0_21 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c21
*+ bl_0_21 br_0_21 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c21
*+ bl_0_21 br_0_21 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c21
*+ bl_0_21 br_0_21 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c21
*+ bl_0_21 br_0_21 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c21
*+ bl_0_21 br_0_21 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c21
*+ bl_0_21 br_0_21 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c21
*+ bl_0_21 br_0_21 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c21
*+ bl_0_21 br_0_21 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c21
*+ bl_0_21 br_0_21 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c21
*+ bl_0_21 br_0_21 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c21
*+ bl_0_21 br_0_21 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c21
*+ bl_0_21 br_0_21 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c21
*+ bl_0_21 br_0_21 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c21
*+ bl_0_21 br_0_21 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c21
*+ bl_0_21 br_0_21 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c21
*+ bl_0_21 br_0_21 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c21
*+ bl_0_21 br_0_21 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c21
*+ bl_0_21 br_0_21 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c21
*+ bl_0_21 br_0_21 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c21
*+ bl_0_21 br_0_21 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c21
*+ bl_0_21 br_0_21 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c21
*+ bl_0_21 br_0_21 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c21
*+ bl_0_21 br_0_21 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c21
*+ bl_0_21 br_0_21 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c21
*+ bl_0_21 br_0_21 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c21
*+ bl_0_21 br_0_21 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c21
*+ bl_0_21 br_0_21 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c21
*+ bl_0_21 br_0_21 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c21
*+ bl_0_21 br_0_21 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c21
*+ bl_0_21 br_0_21 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c21
*+ bl_0_21 br_0_21 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c21
*+ bl_0_21 br_0_21 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c21
*+ bl_0_21 br_0_21 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c21
*+ bl_0_21 br_0_21 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c21
*+ bl_0_21 br_0_21 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c21
*+ bl_0_21 br_0_21 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c21
*+ bl_0_21 br_0_21 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c21
*+ bl_0_21 br_0_21 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c21
*+ bl_0_21 br_0_21 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c21
*+ bl_0_21 br_0_21 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c21
*+ bl_0_21 br_0_21 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c21
*+ bl_0_21 br_0_21 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c21
*+ bl_0_21 br_0_21 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c21
*+ bl_0_21 br_0_21 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c21
*+ bl_0_21 br_0_21 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c21
*+ bl_0_21 br_0_21 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c21
*+ bl_0_21 br_0_21 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c21
*+ bl_0_21 br_0_21 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c21
*+ bl_0_21 br_0_21 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c21
*+ bl_0_21 br_0_21 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c21
*+ bl_0_21 br_0_21 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c21
*+ bl_0_21 br_0_21 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c21
*+ bl_0_21 br_0_21 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c21
*+ bl_0_21 br_0_21 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c21
*+ bl_0_21 br_0_21 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c21
*+ bl_0_21 br_0_21 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c21
*+ bl_0_21 br_0_21 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c21
*+ bl_0_21 br_0_21 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c21
*+ bl_0_21 br_0_21 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c21
*+ bl_0_21 br_0_21 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c21
*+ bl_0_21 br_0_21 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c21
*+ bl_0_21 br_0_21 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c21
*+ bl_0_21 br_0_21 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c21
*+ bl_0_21 br_0_21 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c21
*+ bl_0_21 br_0_21 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c21
*+ bl_0_21 br_0_21 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c21
*+ bl_0_21 br_0_21 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c21
*+ bl_0_21 br_0_21 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c21
*+ bl_0_21 br_0_21 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c21
*+ bl_0_21 br_0_21 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c21
*+ bl_0_21 br_0_21 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c21
*+ bl_0_21 br_0_21 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c21
*+ bl_0_21 br_0_21 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c21
*+ bl_0_21 br_0_21 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c21
*+ bl_0_21 br_0_21 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c21
*+ bl_0_21 br_0_21 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c21
*+ bl_0_21 br_0_21 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c21
*+ bl_0_21 br_0_21 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c21
+ bl_0_21 br_0_21 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c22
+ bl_0_22 br_0_22 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c22
*+ bl_0_22 br_0_22 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c22
*+ bl_0_22 br_0_22 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c22
*+ bl_0_22 br_0_22 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c22
*+ bl_0_22 br_0_22 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c22
*+ bl_0_22 br_0_22 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c22
*+ bl_0_22 br_0_22 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c22
*+ bl_0_22 br_0_22 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c22
*+ bl_0_22 br_0_22 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c22
*+ bl_0_22 br_0_22 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c22
*+ bl_0_22 br_0_22 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c22
*+ bl_0_22 br_0_22 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c22
*+ bl_0_22 br_0_22 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c22
*+ bl_0_22 br_0_22 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c22
*+ bl_0_22 br_0_22 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c22
*+ bl_0_22 br_0_22 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c22
*+ bl_0_22 br_0_22 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c22
*+ bl_0_22 br_0_22 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c22
*+ bl_0_22 br_0_22 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c22
*+ bl_0_22 br_0_22 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c22
*+ bl_0_22 br_0_22 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c22
*+ bl_0_22 br_0_22 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c22
*+ bl_0_22 br_0_22 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c22
*+ bl_0_22 br_0_22 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c22
*+ bl_0_22 br_0_22 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c22
*+ bl_0_22 br_0_22 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c22
*+ bl_0_22 br_0_22 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c22
*+ bl_0_22 br_0_22 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c22
*+ bl_0_22 br_0_22 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c22
*+ bl_0_22 br_0_22 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c22
*+ bl_0_22 br_0_22 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c22
*+ bl_0_22 br_0_22 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c22
*+ bl_0_22 br_0_22 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c22
*+ bl_0_22 br_0_22 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c22
*+ bl_0_22 br_0_22 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c22
*+ bl_0_22 br_0_22 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c22
*+ bl_0_22 br_0_22 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c22
*+ bl_0_22 br_0_22 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c22
*+ bl_0_22 br_0_22 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c22
*+ bl_0_22 br_0_22 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c22
*+ bl_0_22 br_0_22 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c22
*+ bl_0_22 br_0_22 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c22
*+ bl_0_22 br_0_22 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c22
*+ bl_0_22 br_0_22 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c22
*+ bl_0_22 br_0_22 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c22
*+ bl_0_22 br_0_22 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c22
*+ bl_0_22 br_0_22 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c22
*+ bl_0_22 br_0_22 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c22
*+ bl_0_22 br_0_22 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c22
*+ bl_0_22 br_0_22 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c22
*+ bl_0_22 br_0_22 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c22
*+ bl_0_22 br_0_22 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c22
*+ bl_0_22 br_0_22 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c22
*+ bl_0_22 br_0_22 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c22
*+ bl_0_22 br_0_22 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c22
*+ bl_0_22 br_0_22 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c22
*+ bl_0_22 br_0_22 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c22
*+ bl_0_22 br_0_22 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c22
*+ bl_0_22 br_0_22 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c22
*+ bl_0_22 br_0_22 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c22
*+ bl_0_22 br_0_22 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c22
*+ bl_0_22 br_0_22 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c22
*+ bl_0_22 br_0_22 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c22
*+ bl_0_22 br_0_22 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c22
*+ bl_0_22 br_0_22 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c22
*+ bl_0_22 br_0_22 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c22
*+ bl_0_22 br_0_22 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c22
*+ bl_0_22 br_0_22 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c22
*+ bl_0_22 br_0_22 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c22
*+ bl_0_22 br_0_22 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c22
*+ bl_0_22 br_0_22 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c22
*+ bl_0_22 br_0_22 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c22
*+ bl_0_22 br_0_22 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c22
*+ bl_0_22 br_0_22 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c22
*+ bl_0_22 br_0_22 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c22
*+ bl_0_22 br_0_22 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c22
*+ bl_0_22 br_0_22 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c22
*+ bl_0_22 br_0_22 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c22
*+ bl_0_22 br_0_22 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c22
*+ bl_0_22 br_0_22 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c22
*+ bl_0_22 br_0_22 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c22
*+ bl_0_22 br_0_22 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c22
*+ bl_0_22 br_0_22 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c22
*+ bl_0_22 br_0_22 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c22
*+ bl_0_22 br_0_22 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c22
*+ bl_0_22 br_0_22 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c22
*+ bl_0_22 br_0_22 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c22
*+ bl_0_22 br_0_22 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c22
*+ bl_0_22 br_0_22 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c22
*+ bl_0_22 br_0_22 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c22
*+ bl_0_22 br_0_22 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c22
*+ bl_0_22 br_0_22 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c22
*+ bl_0_22 br_0_22 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c22
*+ bl_0_22 br_0_22 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c22
*+ bl_0_22 br_0_22 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c22
*+ bl_0_22 br_0_22 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c22
*+ bl_0_22 br_0_22 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c22
*+ bl_0_22 br_0_22 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c22
*+ bl_0_22 br_0_22 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c22
*+ bl_0_22 br_0_22 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c22
*+ bl_0_22 br_0_22 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c22
*+ bl_0_22 br_0_22 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c22
*+ bl_0_22 br_0_22 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c22
*+ bl_0_22 br_0_22 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c22
*+ bl_0_22 br_0_22 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c22
*+ bl_0_22 br_0_22 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c22
*+ bl_0_22 br_0_22 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c22
*+ bl_0_22 br_0_22 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c22
*+ bl_0_22 br_0_22 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c22
*+ bl_0_22 br_0_22 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c22
*+ bl_0_22 br_0_22 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c22
*+ bl_0_22 br_0_22 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c22
*+ bl_0_22 br_0_22 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c22
*+ bl_0_22 br_0_22 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c22
*+ bl_0_22 br_0_22 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c22
*+ bl_0_22 br_0_22 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c22
*+ bl_0_22 br_0_22 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c22
*+ bl_0_22 br_0_22 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c22
*+ bl_0_22 br_0_22 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c22
*+ bl_0_22 br_0_22 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c22
*+ bl_0_22 br_0_22 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c22
*+ bl_0_22 br_0_22 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c22
*+ bl_0_22 br_0_22 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c22
*+ bl_0_22 br_0_22 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c22
*+ bl_0_22 br_0_22 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c22
*+ bl_0_22 br_0_22 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c22
*+ bl_0_22 br_0_22 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c22
+ bl_0_22 br_0_22 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c23
+ bl_0_23 br_0_23 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c23
*+ bl_0_23 br_0_23 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c23
*+ bl_0_23 br_0_23 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c23
*+ bl_0_23 br_0_23 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c23
*+ bl_0_23 br_0_23 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c23
*+ bl_0_23 br_0_23 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c23
*+ bl_0_23 br_0_23 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c23
*+ bl_0_23 br_0_23 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c23
*+ bl_0_23 br_0_23 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c23
*+ bl_0_23 br_0_23 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c23
*+ bl_0_23 br_0_23 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c23
*+ bl_0_23 br_0_23 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c23
*+ bl_0_23 br_0_23 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c23
*+ bl_0_23 br_0_23 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c23
*+ bl_0_23 br_0_23 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c23
*+ bl_0_23 br_0_23 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c23
*+ bl_0_23 br_0_23 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c23
*+ bl_0_23 br_0_23 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c23
*+ bl_0_23 br_0_23 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c23
*+ bl_0_23 br_0_23 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c23
*+ bl_0_23 br_0_23 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c23
*+ bl_0_23 br_0_23 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c23
*+ bl_0_23 br_0_23 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c23
*+ bl_0_23 br_0_23 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c23
*+ bl_0_23 br_0_23 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c23
*+ bl_0_23 br_0_23 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c23
*+ bl_0_23 br_0_23 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c23
*+ bl_0_23 br_0_23 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c23
*+ bl_0_23 br_0_23 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c23
*+ bl_0_23 br_0_23 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c23
*+ bl_0_23 br_0_23 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c23
*+ bl_0_23 br_0_23 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c23
*+ bl_0_23 br_0_23 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c23
*+ bl_0_23 br_0_23 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c23
*+ bl_0_23 br_0_23 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c23
*+ bl_0_23 br_0_23 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c23
*+ bl_0_23 br_0_23 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c23
*+ bl_0_23 br_0_23 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c23
*+ bl_0_23 br_0_23 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c23
*+ bl_0_23 br_0_23 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c23
*+ bl_0_23 br_0_23 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c23
*+ bl_0_23 br_0_23 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c23
*+ bl_0_23 br_0_23 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c23
*+ bl_0_23 br_0_23 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c23
*+ bl_0_23 br_0_23 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c23
*+ bl_0_23 br_0_23 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c23
*+ bl_0_23 br_0_23 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c23
*+ bl_0_23 br_0_23 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c23
*+ bl_0_23 br_0_23 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c23
*+ bl_0_23 br_0_23 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c23
*+ bl_0_23 br_0_23 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c23
*+ bl_0_23 br_0_23 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c23
*+ bl_0_23 br_0_23 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c23
*+ bl_0_23 br_0_23 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c23
*+ bl_0_23 br_0_23 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c23
*+ bl_0_23 br_0_23 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c23
*+ bl_0_23 br_0_23 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c23
*+ bl_0_23 br_0_23 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c23
*+ bl_0_23 br_0_23 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c23
*+ bl_0_23 br_0_23 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c23
*+ bl_0_23 br_0_23 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c23
*+ bl_0_23 br_0_23 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c23
*+ bl_0_23 br_0_23 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c23
*+ bl_0_23 br_0_23 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c23
*+ bl_0_23 br_0_23 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c23
*+ bl_0_23 br_0_23 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c23
*+ bl_0_23 br_0_23 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c23
*+ bl_0_23 br_0_23 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c23
*+ bl_0_23 br_0_23 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c23
*+ bl_0_23 br_0_23 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c23
*+ bl_0_23 br_0_23 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c23
*+ bl_0_23 br_0_23 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c23
*+ bl_0_23 br_0_23 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c23
*+ bl_0_23 br_0_23 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c23
*+ bl_0_23 br_0_23 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c23
*+ bl_0_23 br_0_23 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c23
*+ bl_0_23 br_0_23 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c23
*+ bl_0_23 br_0_23 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c23
*+ bl_0_23 br_0_23 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c23
*+ bl_0_23 br_0_23 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c23
*+ bl_0_23 br_0_23 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c23
*+ bl_0_23 br_0_23 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c23
*+ bl_0_23 br_0_23 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c23
*+ bl_0_23 br_0_23 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c23
*+ bl_0_23 br_0_23 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c23
*+ bl_0_23 br_0_23 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c23
*+ bl_0_23 br_0_23 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c23
*+ bl_0_23 br_0_23 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c23
*+ bl_0_23 br_0_23 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c23
*+ bl_0_23 br_0_23 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c23
*+ bl_0_23 br_0_23 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c23
*+ bl_0_23 br_0_23 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c23
*+ bl_0_23 br_0_23 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c23
*+ bl_0_23 br_0_23 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c23
*+ bl_0_23 br_0_23 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c23
*+ bl_0_23 br_0_23 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c23
*+ bl_0_23 br_0_23 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c23
*+ bl_0_23 br_0_23 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c23
*+ bl_0_23 br_0_23 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c23
*+ bl_0_23 br_0_23 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c23
*+ bl_0_23 br_0_23 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c23
*+ bl_0_23 br_0_23 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c23
*+ bl_0_23 br_0_23 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c23
*+ bl_0_23 br_0_23 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c23
*+ bl_0_23 br_0_23 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c23
*+ bl_0_23 br_0_23 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c23
*+ bl_0_23 br_0_23 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c23
*+ bl_0_23 br_0_23 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c23
*+ bl_0_23 br_0_23 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c23
*+ bl_0_23 br_0_23 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c23
*+ bl_0_23 br_0_23 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c23
*+ bl_0_23 br_0_23 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c23
*+ bl_0_23 br_0_23 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c23
*+ bl_0_23 br_0_23 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c23
*+ bl_0_23 br_0_23 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c23
*+ bl_0_23 br_0_23 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c23
*+ bl_0_23 br_0_23 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c23
*+ bl_0_23 br_0_23 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c23
*+ bl_0_23 br_0_23 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c23
*+ bl_0_23 br_0_23 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c23
*+ bl_0_23 br_0_23 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c23
*+ bl_0_23 br_0_23 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c23
*+ bl_0_23 br_0_23 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c23
*+ bl_0_23 br_0_23 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c23
*+ bl_0_23 br_0_23 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c23
*+ bl_0_23 br_0_23 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c23
*+ bl_0_23 br_0_23 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c23
+ bl_0_23 br_0_23 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c24
+ bl_0_24 br_0_24 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c24
*+ bl_0_24 br_0_24 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c24
*+ bl_0_24 br_0_24 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c24
*+ bl_0_24 br_0_24 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c24
*+ bl_0_24 br_0_24 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c24
*+ bl_0_24 br_0_24 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c24
*+ bl_0_24 br_0_24 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c24
*+ bl_0_24 br_0_24 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c24
*+ bl_0_24 br_0_24 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c24
*+ bl_0_24 br_0_24 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c24
*+ bl_0_24 br_0_24 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c24
*+ bl_0_24 br_0_24 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c24
*+ bl_0_24 br_0_24 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c24
*+ bl_0_24 br_0_24 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c24
*+ bl_0_24 br_0_24 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c24
*+ bl_0_24 br_0_24 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c24
*+ bl_0_24 br_0_24 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c24
*+ bl_0_24 br_0_24 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c24
*+ bl_0_24 br_0_24 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c24
*+ bl_0_24 br_0_24 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c24
*+ bl_0_24 br_0_24 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c24
*+ bl_0_24 br_0_24 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c24
*+ bl_0_24 br_0_24 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c24
*+ bl_0_24 br_0_24 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c24
*+ bl_0_24 br_0_24 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c24
*+ bl_0_24 br_0_24 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c24
*+ bl_0_24 br_0_24 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c24
*+ bl_0_24 br_0_24 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c24
*+ bl_0_24 br_0_24 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c24
*+ bl_0_24 br_0_24 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c24
*+ bl_0_24 br_0_24 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c24
*+ bl_0_24 br_0_24 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c24
*+ bl_0_24 br_0_24 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c24
*+ bl_0_24 br_0_24 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c24
*+ bl_0_24 br_0_24 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c24
*+ bl_0_24 br_0_24 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c24
*+ bl_0_24 br_0_24 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c24
*+ bl_0_24 br_0_24 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c24
*+ bl_0_24 br_0_24 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c24
*+ bl_0_24 br_0_24 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c24
*+ bl_0_24 br_0_24 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c24
*+ bl_0_24 br_0_24 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c24
*+ bl_0_24 br_0_24 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c24
*+ bl_0_24 br_0_24 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c24
*+ bl_0_24 br_0_24 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c24
*+ bl_0_24 br_0_24 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c24
*+ bl_0_24 br_0_24 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c24
*+ bl_0_24 br_0_24 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c24
*+ bl_0_24 br_0_24 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c24
*+ bl_0_24 br_0_24 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c24
*+ bl_0_24 br_0_24 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c24
*+ bl_0_24 br_0_24 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c24
*+ bl_0_24 br_0_24 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c24
*+ bl_0_24 br_0_24 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c24
*+ bl_0_24 br_0_24 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c24
*+ bl_0_24 br_0_24 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c24
*+ bl_0_24 br_0_24 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c24
*+ bl_0_24 br_0_24 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c24
*+ bl_0_24 br_0_24 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c24
*+ bl_0_24 br_0_24 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c24
*+ bl_0_24 br_0_24 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c24
*+ bl_0_24 br_0_24 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c24
*+ bl_0_24 br_0_24 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c24
*+ bl_0_24 br_0_24 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c24
*+ bl_0_24 br_0_24 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c24
*+ bl_0_24 br_0_24 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c24
*+ bl_0_24 br_0_24 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c24
*+ bl_0_24 br_0_24 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c24
*+ bl_0_24 br_0_24 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c24
*+ bl_0_24 br_0_24 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c24
*+ bl_0_24 br_0_24 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c24
*+ bl_0_24 br_0_24 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c24
*+ bl_0_24 br_0_24 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c24
*+ bl_0_24 br_0_24 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c24
*+ bl_0_24 br_0_24 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c24
*+ bl_0_24 br_0_24 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c24
*+ bl_0_24 br_0_24 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c24
*+ bl_0_24 br_0_24 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c24
*+ bl_0_24 br_0_24 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c24
*+ bl_0_24 br_0_24 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c24
*+ bl_0_24 br_0_24 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c24
*+ bl_0_24 br_0_24 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c24
*+ bl_0_24 br_0_24 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c24
*+ bl_0_24 br_0_24 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c24
*+ bl_0_24 br_0_24 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c24
*+ bl_0_24 br_0_24 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c24
*+ bl_0_24 br_0_24 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c24
*+ bl_0_24 br_0_24 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c24
*+ bl_0_24 br_0_24 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c24
*+ bl_0_24 br_0_24 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c24
*+ bl_0_24 br_0_24 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c24
*+ bl_0_24 br_0_24 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c24
*+ bl_0_24 br_0_24 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c24
*+ bl_0_24 br_0_24 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c24
*+ bl_0_24 br_0_24 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c24
*+ bl_0_24 br_0_24 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c24
*+ bl_0_24 br_0_24 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c24
*+ bl_0_24 br_0_24 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c24
*+ bl_0_24 br_0_24 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c24
*+ bl_0_24 br_0_24 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c24
*+ bl_0_24 br_0_24 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c24
*+ bl_0_24 br_0_24 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c24
*+ bl_0_24 br_0_24 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c24
*+ bl_0_24 br_0_24 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c24
*+ bl_0_24 br_0_24 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c24
*+ bl_0_24 br_0_24 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c24
*+ bl_0_24 br_0_24 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c24
*+ bl_0_24 br_0_24 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c24
*+ bl_0_24 br_0_24 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c24
*+ bl_0_24 br_0_24 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c24
*+ bl_0_24 br_0_24 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c24
*+ bl_0_24 br_0_24 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c24
*+ bl_0_24 br_0_24 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c24
*+ bl_0_24 br_0_24 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c24
*+ bl_0_24 br_0_24 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c24
*+ bl_0_24 br_0_24 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c24
*+ bl_0_24 br_0_24 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c24
*+ bl_0_24 br_0_24 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c24
*+ bl_0_24 br_0_24 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c24
*+ bl_0_24 br_0_24 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c24
*+ bl_0_24 br_0_24 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c24
*+ bl_0_24 br_0_24 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c24
*+ bl_0_24 br_0_24 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c24
*+ bl_0_24 br_0_24 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c24
*+ bl_0_24 br_0_24 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c24
*+ bl_0_24 br_0_24 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c24
*+ bl_0_24 br_0_24 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c24
+ bl_0_24 br_0_24 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c25
+ bl_0_25 br_0_25 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c25
*+ bl_0_25 br_0_25 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c25
*+ bl_0_25 br_0_25 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c25
*+ bl_0_25 br_0_25 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c25
*+ bl_0_25 br_0_25 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c25
*+ bl_0_25 br_0_25 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c25
*+ bl_0_25 br_0_25 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c25
*+ bl_0_25 br_0_25 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c25
*+ bl_0_25 br_0_25 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c25
*+ bl_0_25 br_0_25 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c25
*+ bl_0_25 br_0_25 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c25
*+ bl_0_25 br_0_25 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c25
*+ bl_0_25 br_0_25 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c25
*+ bl_0_25 br_0_25 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c25
*+ bl_0_25 br_0_25 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c25
*+ bl_0_25 br_0_25 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c25
*+ bl_0_25 br_0_25 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c25
*+ bl_0_25 br_0_25 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c25
*+ bl_0_25 br_0_25 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c25
*+ bl_0_25 br_0_25 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c25
*+ bl_0_25 br_0_25 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c25
*+ bl_0_25 br_0_25 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c25
*+ bl_0_25 br_0_25 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c25
*+ bl_0_25 br_0_25 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c25
*+ bl_0_25 br_0_25 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c25
*+ bl_0_25 br_0_25 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c25
*+ bl_0_25 br_0_25 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c25
*+ bl_0_25 br_0_25 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c25
*+ bl_0_25 br_0_25 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c25
*+ bl_0_25 br_0_25 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c25
*+ bl_0_25 br_0_25 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c25
*+ bl_0_25 br_0_25 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c25
*+ bl_0_25 br_0_25 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c25
*+ bl_0_25 br_0_25 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c25
*+ bl_0_25 br_0_25 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c25
*+ bl_0_25 br_0_25 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c25
*+ bl_0_25 br_0_25 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c25
*+ bl_0_25 br_0_25 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c25
*+ bl_0_25 br_0_25 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c25
*+ bl_0_25 br_0_25 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c25
*+ bl_0_25 br_0_25 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c25
*+ bl_0_25 br_0_25 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c25
*+ bl_0_25 br_0_25 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c25
*+ bl_0_25 br_0_25 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c25
*+ bl_0_25 br_0_25 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c25
*+ bl_0_25 br_0_25 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c25
*+ bl_0_25 br_0_25 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c25
*+ bl_0_25 br_0_25 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c25
*+ bl_0_25 br_0_25 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c25
*+ bl_0_25 br_0_25 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c25
*+ bl_0_25 br_0_25 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c25
*+ bl_0_25 br_0_25 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c25
*+ bl_0_25 br_0_25 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c25
*+ bl_0_25 br_0_25 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c25
*+ bl_0_25 br_0_25 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c25
*+ bl_0_25 br_0_25 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c25
*+ bl_0_25 br_0_25 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c25
*+ bl_0_25 br_0_25 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c25
*+ bl_0_25 br_0_25 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c25
*+ bl_0_25 br_0_25 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c25
*+ bl_0_25 br_0_25 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c25
*+ bl_0_25 br_0_25 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c25
*+ bl_0_25 br_0_25 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c25
*+ bl_0_25 br_0_25 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c25
*+ bl_0_25 br_0_25 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c25
*+ bl_0_25 br_0_25 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c25
*+ bl_0_25 br_0_25 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c25
*+ bl_0_25 br_0_25 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c25
*+ bl_0_25 br_0_25 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c25
*+ bl_0_25 br_0_25 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c25
*+ bl_0_25 br_0_25 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c25
*+ bl_0_25 br_0_25 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c25
*+ bl_0_25 br_0_25 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c25
*+ bl_0_25 br_0_25 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c25
*+ bl_0_25 br_0_25 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c25
*+ bl_0_25 br_0_25 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c25
*+ bl_0_25 br_0_25 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c25
*+ bl_0_25 br_0_25 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c25
*+ bl_0_25 br_0_25 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c25
*+ bl_0_25 br_0_25 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c25
*+ bl_0_25 br_0_25 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c25
*+ bl_0_25 br_0_25 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c25
*+ bl_0_25 br_0_25 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c25
*+ bl_0_25 br_0_25 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c25
*+ bl_0_25 br_0_25 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c25
*+ bl_0_25 br_0_25 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c25
*+ bl_0_25 br_0_25 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c25
*+ bl_0_25 br_0_25 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c25
*+ bl_0_25 br_0_25 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c25
*+ bl_0_25 br_0_25 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c25
*+ bl_0_25 br_0_25 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c25
*+ bl_0_25 br_0_25 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c25
*+ bl_0_25 br_0_25 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c25
*+ bl_0_25 br_0_25 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c25
*+ bl_0_25 br_0_25 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c25
*+ bl_0_25 br_0_25 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c25
*+ bl_0_25 br_0_25 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c25
*+ bl_0_25 br_0_25 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c25
*+ bl_0_25 br_0_25 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c25
*+ bl_0_25 br_0_25 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c25
*+ bl_0_25 br_0_25 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c25
*+ bl_0_25 br_0_25 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c25
*+ bl_0_25 br_0_25 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c25
*+ bl_0_25 br_0_25 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c25
*+ bl_0_25 br_0_25 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c25
*+ bl_0_25 br_0_25 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c25
*+ bl_0_25 br_0_25 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c25
*+ bl_0_25 br_0_25 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c25
*+ bl_0_25 br_0_25 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c25
*+ bl_0_25 br_0_25 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c25
*+ bl_0_25 br_0_25 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c25
*+ bl_0_25 br_0_25 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c25
*+ bl_0_25 br_0_25 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c25
*+ bl_0_25 br_0_25 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c25
*+ bl_0_25 br_0_25 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c25
*+ bl_0_25 br_0_25 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c25
*+ bl_0_25 br_0_25 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c25
*+ bl_0_25 br_0_25 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c25
*+ bl_0_25 br_0_25 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c25
*+ bl_0_25 br_0_25 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c25
*+ bl_0_25 br_0_25 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c25
*+ bl_0_25 br_0_25 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c25
*+ bl_0_25 br_0_25 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c25
*+ bl_0_25 br_0_25 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c25
*+ bl_0_25 br_0_25 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c25
*+ bl_0_25 br_0_25 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c25
*+ bl_0_25 br_0_25 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c25
+ bl_0_25 br_0_25 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c26
+ bl_0_26 br_0_26 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c26
*+ bl_0_26 br_0_26 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c26
*+ bl_0_26 br_0_26 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c26
*+ bl_0_26 br_0_26 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c26
*+ bl_0_26 br_0_26 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c26
*+ bl_0_26 br_0_26 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c26
*+ bl_0_26 br_0_26 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c26
*+ bl_0_26 br_0_26 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c26
*+ bl_0_26 br_0_26 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c26
*+ bl_0_26 br_0_26 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c26
*+ bl_0_26 br_0_26 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c26
*+ bl_0_26 br_0_26 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c26
*+ bl_0_26 br_0_26 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c26
*+ bl_0_26 br_0_26 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c26
*+ bl_0_26 br_0_26 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c26
*+ bl_0_26 br_0_26 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c26
*+ bl_0_26 br_0_26 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c26
*+ bl_0_26 br_0_26 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c26
*+ bl_0_26 br_0_26 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c26
*+ bl_0_26 br_0_26 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c26
*+ bl_0_26 br_0_26 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c26
*+ bl_0_26 br_0_26 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c26
*+ bl_0_26 br_0_26 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c26
*+ bl_0_26 br_0_26 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c26
*+ bl_0_26 br_0_26 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c26
*+ bl_0_26 br_0_26 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c26
*+ bl_0_26 br_0_26 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c26
*+ bl_0_26 br_0_26 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c26
*+ bl_0_26 br_0_26 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c26
*+ bl_0_26 br_0_26 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c26
*+ bl_0_26 br_0_26 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c26
*+ bl_0_26 br_0_26 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c26
*+ bl_0_26 br_0_26 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c26
*+ bl_0_26 br_0_26 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c26
*+ bl_0_26 br_0_26 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c26
*+ bl_0_26 br_0_26 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c26
*+ bl_0_26 br_0_26 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c26
*+ bl_0_26 br_0_26 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c26
*+ bl_0_26 br_0_26 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c26
*+ bl_0_26 br_0_26 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c26
*+ bl_0_26 br_0_26 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c26
*+ bl_0_26 br_0_26 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c26
*+ bl_0_26 br_0_26 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c26
*+ bl_0_26 br_0_26 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c26
*+ bl_0_26 br_0_26 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c26
*+ bl_0_26 br_0_26 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c26
*+ bl_0_26 br_0_26 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c26
*+ bl_0_26 br_0_26 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c26
*+ bl_0_26 br_0_26 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c26
*+ bl_0_26 br_0_26 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c26
*+ bl_0_26 br_0_26 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c26
*+ bl_0_26 br_0_26 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c26
*+ bl_0_26 br_0_26 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c26
*+ bl_0_26 br_0_26 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c26
*+ bl_0_26 br_0_26 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c26
*+ bl_0_26 br_0_26 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c26
*+ bl_0_26 br_0_26 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c26
*+ bl_0_26 br_0_26 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c26
*+ bl_0_26 br_0_26 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c26
*+ bl_0_26 br_0_26 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c26
*+ bl_0_26 br_0_26 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c26
*+ bl_0_26 br_0_26 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c26
*+ bl_0_26 br_0_26 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c26
*+ bl_0_26 br_0_26 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c26
*+ bl_0_26 br_0_26 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c26
*+ bl_0_26 br_0_26 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c26
*+ bl_0_26 br_0_26 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c26
*+ bl_0_26 br_0_26 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c26
*+ bl_0_26 br_0_26 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c26
*+ bl_0_26 br_0_26 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c26
*+ bl_0_26 br_0_26 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c26
*+ bl_0_26 br_0_26 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c26
*+ bl_0_26 br_0_26 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c26
*+ bl_0_26 br_0_26 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c26
*+ bl_0_26 br_0_26 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c26
*+ bl_0_26 br_0_26 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c26
*+ bl_0_26 br_0_26 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c26
*+ bl_0_26 br_0_26 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c26
*+ bl_0_26 br_0_26 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c26
*+ bl_0_26 br_0_26 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c26
*+ bl_0_26 br_0_26 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c26
*+ bl_0_26 br_0_26 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c26
*+ bl_0_26 br_0_26 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c26
*+ bl_0_26 br_0_26 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c26
*+ bl_0_26 br_0_26 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c26
*+ bl_0_26 br_0_26 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c26
*+ bl_0_26 br_0_26 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c26
*+ bl_0_26 br_0_26 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c26
*+ bl_0_26 br_0_26 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c26
*+ bl_0_26 br_0_26 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c26
*+ bl_0_26 br_0_26 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c26
*+ bl_0_26 br_0_26 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c26
*+ bl_0_26 br_0_26 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c26
*+ bl_0_26 br_0_26 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c26
*+ bl_0_26 br_0_26 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c26
*+ bl_0_26 br_0_26 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c26
*+ bl_0_26 br_0_26 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c26
*+ bl_0_26 br_0_26 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c26
*+ bl_0_26 br_0_26 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c26
*+ bl_0_26 br_0_26 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c26
*+ bl_0_26 br_0_26 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c26
*+ bl_0_26 br_0_26 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c26
*+ bl_0_26 br_0_26 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c26
*+ bl_0_26 br_0_26 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c26
*+ bl_0_26 br_0_26 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c26
*+ bl_0_26 br_0_26 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c26
*+ bl_0_26 br_0_26 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c26
*+ bl_0_26 br_0_26 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c26
*+ bl_0_26 br_0_26 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c26
*+ bl_0_26 br_0_26 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c26
*+ bl_0_26 br_0_26 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c26
*+ bl_0_26 br_0_26 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c26
*+ bl_0_26 br_0_26 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c26
*+ bl_0_26 br_0_26 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c26
*+ bl_0_26 br_0_26 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c26
*+ bl_0_26 br_0_26 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c26
*+ bl_0_26 br_0_26 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c26
*+ bl_0_26 br_0_26 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c26
*+ bl_0_26 br_0_26 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c26
*+ bl_0_26 br_0_26 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c26
*+ bl_0_26 br_0_26 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c26
*+ bl_0_26 br_0_26 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c26
*+ bl_0_26 br_0_26 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c26
*+ bl_0_26 br_0_26 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c26
*+ bl_0_26 br_0_26 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c26
*+ bl_0_26 br_0_26 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c26
*+ bl_0_26 br_0_26 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c26
+ bl_0_26 br_0_26 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c27
+ bl_0_27 br_0_27 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c27
*+ bl_0_27 br_0_27 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c27
*+ bl_0_27 br_0_27 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c27
*+ bl_0_27 br_0_27 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c27
*+ bl_0_27 br_0_27 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c27
*+ bl_0_27 br_0_27 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c27
*+ bl_0_27 br_0_27 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c27
*+ bl_0_27 br_0_27 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c27
*+ bl_0_27 br_0_27 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c27
*+ bl_0_27 br_0_27 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c27
*+ bl_0_27 br_0_27 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c27
*+ bl_0_27 br_0_27 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c27
*+ bl_0_27 br_0_27 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c27
*+ bl_0_27 br_0_27 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c27
*+ bl_0_27 br_0_27 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c27
*+ bl_0_27 br_0_27 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c27
*+ bl_0_27 br_0_27 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c27
*+ bl_0_27 br_0_27 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c27
*+ bl_0_27 br_0_27 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c27
*+ bl_0_27 br_0_27 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c27
*+ bl_0_27 br_0_27 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c27
*+ bl_0_27 br_0_27 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c27
*+ bl_0_27 br_0_27 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c27
*+ bl_0_27 br_0_27 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c27
*+ bl_0_27 br_0_27 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c27
*+ bl_0_27 br_0_27 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c27
*+ bl_0_27 br_0_27 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c27
*+ bl_0_27 br_0_27 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c27
*+ bl_0_27 br_0_27 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c27
*+ bl_0_27 br_0_27 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c27
*+ bl_0_27 br_0_27 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c27
*+ bl_0_27 br_0_27 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c27
*+ bl_0_27 br_0_27 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c27
*+ bl_0_27 br_0_27 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c27
*+ bl_0_27 br_0_27 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c27
*+ bl_0_27 br_0_27 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c27
*+ bl_0_27 br_0_27 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c27
*+ bl_0_27 br_0_27 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c27
*+ bl_0_27 br_0_27 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c27
*+ bl_0_27 br_0_27 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c27
*+ bl_0_27 br_0_27 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c27
*+ bl_0_27 br_0_27 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c27
*+ bl_0_27 br_0_27 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c27
*+ bl_0_27 br_0_27 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c27
*+ bl_0_27 br_0_27 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c27
*+ bl_0_27 br_0_27 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c27
*+ bl_0_27 br_0_27 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c27
*+ bl_0_27 br_0_27 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c27
*+ bl_0_27 br_0_27 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c27
*+ bl_0_27 br_0_27 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c27
*+ bl_0_27 br_0_27 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c27
*+ bl_0_27 br_0_27 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c27
*+ bl_0_27 br_0_27 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c27
*+ bl_0_27 br_0_27 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c27
*+ bl_0_27 br_0_27 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c27
*+ bl_0_27 br_0_27 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c27
*+ bl_0_27 br_0_27 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c27
*+ bl_0_27 br_0_27 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c27
*+ bl_0_27 br_0_27 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c27
*+ bl_0_27 br_0_27 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c27
*+ bl_0_27 br_0_27 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c27
*+ bl_0_27 br_0_27 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c27
*+ bl_0_27 br_0_27 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c27
*+ bl_0_27 br_0_27 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c27
*+ bl_0_27 br_0_27 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c27
*+ bl_0_27 br_0_27 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c27
*+ bl_0_27 br_0_27 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c27
*+ bl_0_27 br_0_27 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c27
*+ bl_0_27 br_0_27 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c27
*+ bl_0_27 br_0_27 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c27
*+ bl_0_27 br_0_27 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c27
*+ bl_0_27 br_0_27 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c27
*+ bl_0_27 br_0_27 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c27
*+ bl_0_27 br_0_27 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c27
*+ bl_0_27 br_0_27 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c27
*+ bl_0_27 br_0_27 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c27
*+ bl_0_27 br_0_27 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c27
*+ bl_0_27 br_0_27 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c27
*+ bl_0_27 br_0_27 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c27
*+ bl_0_27 br_0_27 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c27
*+ bl_0_27 br_0_27 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c27
*+ bl_0_27 br_0_27 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c27
*+ bl_0_27 br_0_27 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c27
*+ bl_0_27 br_0_27 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c27
*+ bl_0_27 br_0_27 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c27
*+ bl_0_27 br_0_27 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c27
*+ bl_0_27 br_0_27 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c27
*+ bl_0_27 br_0_27 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c27
*+ bl_0_27 br_0_27 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c27
*+ bl_0_27 br_0_27 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c27
*+ bl_0_27 br_0_27 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c27
*+ bl_0_27 br_0_27 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c27
*+ bl_0_27 br_0_27 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c27
*+ bl_0_27 br_0_27 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c27
*+ bl_0_27 br_0_27 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c27
*+ bl_0_27 br_0_27 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c27
*+ bl_0_27 br_0_27 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c27
*+ bl_0_27 br_0_27 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c27
*+ bl_0_27 br_0_27 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c27
*+ bl_0_27 br_0_27 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c27
*+ bl_0_27 br_0_27 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c27
*+ bl_0_27 br_0_27 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c27
*+ bl_0_27 br_0_27 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c27
*+ bl_0_27 br_0_27 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c27
*+ bl_0_27 br_0_27 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c27
*+ bl_0_27 br_0_27 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c27
*+ bl_0_27 br_0_27 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c27
*+ bl_0_27 br_0_27 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c27
*+ bl_0_27 br_0_27 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c27
*+ bl_0_27 br_0_27 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c27
*+ bl_0_27 br_0_27 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c27
*+ bl_0_27 br_0_27 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c27
*+ bl_0_27 br_0_27 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c27
*+ bl_0_27 br_0_27 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c27
*+ bl_0_27 br_0_27 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c27
*+ bl_0_27 br_0_27 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c27
*+ bl_0_27 br_0_27 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c27
*+ bl_0_27 br_0_27 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c27
*+ bl_0_27 br_0_27 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c27
*+ bl_0_27 br_0_27 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c27
*+ bl_0_27 br_0_27 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c27
*+ bl_0_27 br_0_27 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c27
*+ bl_0_27 br_0_27 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c27
*+ bl_0_27 br_0_27 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c27
*+ bl_0_27 br_0_27 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c27
*+ bl_0_27 br_0_27 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c27
*+ bl_0_27 br_0_27 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c27
+ bl_0_27 br_0_27 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c28
+ bl_0_28 br_0_28 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c28
*+ bl_0_28 br_0_28 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c28
*+ bl_0_28 br_0_28 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c28
*+ bl_0_28 br_0_28 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c28
*+ bl_0_28 br_0_28 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c28
*+ bl_0_28 br_0_28 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c28
*+ bl_0_28 br_0_28 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c28
*+ bl_0_28 br_0_28 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c28
*+ bl_0_28 br_0_28 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c28
*+ bl_0_28 br_0_28 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c28
*+ bl_0_28 br_0_28 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c28
*+ bl_0_28 br_0_28 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c28
*+ bl_0_28 br_0_28 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c28
*+ bl_0_28 br_0_28 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c28
*+ bl_0_28 br_0_28 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c28
*+ bl_0_28 br_0_28 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c28
*+ bl_0_28 br_0_28 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c28
*+ bl_0_28 br_0_28 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c28
*+ bl_0_28 br_0_28 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c28
*+ bl_0_28 br_0_28 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c28
*+ bl_0_28 br_0_28 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c28
*+ bl_0_28 br_0_28 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c28
*+ bl_0_28 br_0_28 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c28
*+ bl_0_28 br_0_28 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c28
*+ bl_0_28 br_0_28 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c28
*+ bl_0_28 br_0_28 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c28
*+ bl_0_28 br_0_28 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c28
*+ bl_0_28 br_0_28 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c28
*+ bl_0_28 br_0_28 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c28
*+ bl_0_28 br_0_28 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c28
*+ bl_0_28 br_0_28 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c28
*+ bl_0_28 br_0_28 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c28
*+ bl_0_28 br_0_28 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c28
*+ bl_0_28 br_0_28 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c28
*+ bl_0_28 br_0_28 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c28
*+ bl_0_28 br_0_28 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c28
*+ bl_0_28 br_0_28 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c28
*+ bl_0_28 br_0_28 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c28
*+ bl_0_28 br_0_28 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c28
*+ bl_0_28 br_0_28 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c28
*+ bl_0_28 br_0_28 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c28
*+ bl_0_28 br_0_28 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c28
*+ bl_0_28 br_0_28 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c28
*+ bl_0_28 br_0_28 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c28
*+ bl_0_28 br_0_28 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c28
*+ bl_0_28 br_0_28 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c28
*+ bl_0_28 br_0_28 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c28
*+ bl_0_28 br_0_28 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c28
*+ bl_0_28 br_0_28 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c28
*+ bl_0_28 br_0_28 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c28
*+ bl_0_28 br_0_28 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c28
*+ bl_0_28 br_0_28 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c28
*+ bl_0_28 br_0_28 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c28
*+ bl_0_28 br_0_28 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c28
*+ bl_0_28 br_0_28 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c28
*+ bl_0_28 br_0_28 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c28
*+ bl_0_28 br_0_28 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c28
*+ bl_0_28 br_0_28 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c28
*+ bl_0_28 br_0_28 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c28
*+ bl_0_28 br_0_28 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c28
*+ bl_0_28 br_0_28 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c28
*+ bl_0_28 br_0_28 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c28
*+ bl_0_28 br_0_28 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c28
*+ bl_0_28 br_0_28 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c28
*+ bl_0_28 br_0_28 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c28
*+ bl_0_28 br_0_28 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c28
*+ bl_0_28 br_0_28 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c28
*+ bl_0_28 br_0_28 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c28
*+ bl_0_28 br_0_28 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c28
*+ bl_0_28 br_0_28 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c28
*+ bl_0_28 br_0_28 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c28
*+ bl_0_28 br_0_28 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c28
*+ bl_0_28 br_0_28 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c28
*+ bl_0_28 br_0_28 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c28
*+ bl_0_28 br_0_28 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c28
*+ bl_0_28 br_0_28 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c28
*+ bl_0_28 br_0_28 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c28
*+ bl_0_28 br_0_28 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c28
*+ bl_0_28 br_0_28 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c28
*+ bl_0_28 br_0_28 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c28
*+ bl_0_28 br_0_28 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c28
*+ bl_0_28 br_0_28 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c28
*+ bl_0_28 br_0_28 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c28
*+ bl_0_28 br_0_28 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c28
*+ bl_0_28 br_0_28 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c28
*+ bl_0_28 br_0_28 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c28
*+ bl_0_28 br_0_28 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c28
*+ bl_0_28 br_0_28 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c28
*+ bl_0_28 br_0_28 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c28
*+ bl_0_28 br_0_28 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c28
*+ bl_0_28 br_0_28 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c28
*+ bl_0_28 br_0_28 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c28
*+ bl_0_28 br_0_28 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c28
*+ bl_0_28 br_0_28 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c28
*+ bl_0_28 br_0_28 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c28
*+ bl_0_28 br_0_28 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c28
*+ bl_0_28 br_0_28 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c28
*+ bl_0_28 br_0_28 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c28
*+ bl_0_28 br_0_28 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c28
*+ bl_0_28 br_0_28 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c28
*+ bl_0_28 br_0_28 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c28
*+ bl_0_28 br_0_28 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c28
*+ bl_0_28 br_0_28 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c28
*+ bl_0_28 br_0_28 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c28
*+ bl_0_28 br_0_28 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c28
*+ bl_0_28 br_0_28 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c28
*+ bl_0_28 br_0_28 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c28
*+ bl_0_28 br_0_28 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c28
*+ bl_0_28 br_0_28 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c28
*+ bl_0_28 br_0_28 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c28
*+ bl_0_28 br_0_28 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c28
*+ bl_0_28 br_0_28 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c28
*+ bl_0_28 br_0_28 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c28
*+ bl_0_28 br_0_28 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c28
*+ bl_0_28 br_0_28 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c28
*+ bl_0_28 br_0_28 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c28
*+ bl_0_28 br_0_28 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c28
*+ bl_0_28 br_0_28 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c28
*+ bl_0_28 br_0_28 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c28
*+ bl_0_28 br_0_28 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c28
*+ bl_0_28 br_0_28 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c28
*+ bl_0_28 br_0_28 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c28
*+ bl_0_28 br_0_28 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c28
*+ bl_0_28 br_0_28 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c28
*+ bl_0_28 br_0_28 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c28
*+ bl_0_28 br_0_28 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c28
*+ bl_0_28 br_0_28 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c28
+ bl_0_28 br_0_28 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c29
+ bl_0_29 br_0_29 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c29
*+ bl_0_29 br_0_29 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c29
*+ bl_0_29 br_0_29 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c29
*+ bl_0_29 br_0_29 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c29
*+ bl_0_29 br_0_29 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c29
*+ bl_0_29 br_0_29 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c29
*+ bl_0_29 br_0_29 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c29
*+ bl_0_29 br_0_29 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c29
*+ bl_0_29 br_0_29 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c29
*+ bl_0_29 br_0_29 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c29
*+ bl_0_29 br_0_29 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c29
*+ bl_0_29 br_0_29 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c29
*+ bl_0_29 br_0_29 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c29
*+ bl_0_29 br_0_29 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c29
*+ bl_0_29 br_0_29 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c29
*+ bl_0_29 br_0_29 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c29
*+ bl_0_29 br_0_29 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c29
*+ bl_0_29 br_0_29 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c29
*+ bl_0_29 br_0_29 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c29
*+ bl_0_29 br_0_29 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c29
*+ bl_0_29 br_0_29 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c29
*+ bl_0_29 br_0_29 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c29
*+ bl_0_29 br_0_29 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c29
*+ bl_0_29 br_0_29 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c29
*+ bl_0_29 br_0_29 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c29
*+ bl_0_29 br_0_29 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c29
*+ bl_0_29 br_0_29 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c29
*+ bl_0_29 br_0_29 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c29
*+ bl_0_29 br_0_29 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c29
*+ bl_0_29 br_0_29 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c29
*+ bl_0_29 br_0_29 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c29
*+ bl_0_29 br_0_29 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c29
*+ bl_0_29 br_0_29 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c29
*+ bl_0_29 br_0_29 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c29
*+ bl_0_29 br_0_29 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c29
*+ bl_0_29 br_0_29 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c29
*+ bl_0_29 br_0_29 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c29
*+ bl_0_29 br_0_29 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c29
*+ bl_0_29 br_0_29 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c29
*+ bl_0_29 br_0_29 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c29
*+ bl_0_29 br_0_29 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c29
*+ bl_0_29 br_0_29 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c29
*+ bl_0_29 br_0_29 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c29
*+ bl_0_29 br_0_29 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c29
*+ bl_0_29 br_0_29 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c29
*+ bl_0_29 br_0_29 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c29
*+ bl_0_29 br_0_29 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c29
*+ bl_0_29 br_0_29 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c29
*+ bl_0_29 br_0_29 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c29
*+ bl_0_29 br_0_29 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c29
*+ bl_0_29 br_0_29 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c29
*+ bl_0_29 br_0_29 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c29
*+ bl_0_29 br_0_29 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c29
*+ bl_0_29 br_0_29 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c29
*+ bl_0_29 br_0_29 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c29
*+ bl_0_29 br_0_29 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c29
*+ bl_0_29 br_0_29 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c29
*+ bl_0_29 br_0_29 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c29
*+ bl_0_29 br_0_29 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c29
*+ bl_0_29 br_0_29 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c29
*+ bl_0_29 br_0_29 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c29
*+ bl_0_29 br_0_29 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c29
*+ bl_0_29 br_0_29 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c29
*+ bl_0_29 br_0_29 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c29
*+ bl_0_29 br_0_29 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c29
*+ bl_0_29 br_0_29 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c29
*+ bl_0_29 br_0_29 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c29
*+ bl_0_29 br_0_29 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c29
*+ bl_0_29 br_0_29 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c29
*+ bl_0_29 br_0_29 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c29
*+ bl_0_29 br_0_29 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c29
*+ bl_0_29 br_0_29 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c29
*+ bl_0_29 br_0_29 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c29
*+ bl_0_29 br_0_29 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c29
*+ bl_0_29 br_0_29 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c29
*+ bl_0_29 br_0_29 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c29
*+ bl_0_29 br_0_29 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c29
*+ bl_0_29 br_0_29 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c29
*+ bl_0_29 br_0_29 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c29
*+ bl_0_29 br_0_29 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c29
*+ bl_0_29 br_0_29 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c29
*+ bl_0_29 br_0_29 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c29
*+ bl_0_29 br_0_29 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c29
*+ bl_0_29 br_0_29 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c29
*+ bl_0_29 br_0_29 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c29
*+ bl_0_29 br_0_29 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c29
*+ bl_0_29 br_0_29 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c29
*+ bl_0_29 br_0_29 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c29
*+ bl_0_29 br_0_29 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c29
*+ bl_0_29 br_0_29 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c29
*+ bl_0_29 br_0_29 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c29
*+ bl_0_29 br_0_29 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c29
*+ bl_0_29 br_0_29 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c29
*+ bl_0_29 br_0_29 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c29
*+ bl_0_29 br_0_29 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c29
*+ bl_0_29 br_0_29 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c29
*+ bl_0_29 br_0_29 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c29
*+ bl_0_29 br_0_29 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c29
*+ bl_0_29 br_0_29 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c29
*+ bl_0_29 br_0_29 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c29
*+ bl_0_29 br_0_29 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c29
*+ bl_0_29 br_0_29 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c29
*+ bl_0_29 br_0_29 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c29
*+ bl_0_29 br_0_29 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c29
*+ bl_0_29 br_0_29 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c29
*+ bl_0_29 br_0_29 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c29
*+ bl_0_29 br_0_29 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c29
*+ bl_0_29 br_0_29 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c29
*+ bl_0_29 br_0_29 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c29
*+ bl_0_29 br_0_29 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c29
*+ bl_0_29 br_0_29 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c29
*+ bl_0_29 br_0_29 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c29
*+ bl_0_29 br_0_29 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c29
*+ bl_0_29 br_0_29 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c29
*+ bl_0_29 br_0_29 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c29
*+ bl_0_29 br_0_29 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c29
*+ bl_0_29 br_0_29 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c29
*+ bl_0_29 br_0_29 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c29
*+ bl_0_29 br_0_29 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c29
*+ bl_0_29 br_0_29 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c29
*+ bl_0_29 br_0_29 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c29
*+ bl_0_29 br_0_29 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c29
*+ bl_0_29 br_0_29 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c29
*+ bl_0_29 br_0_29 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c29
*+ bl_0_29 br_0_29 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c29
*+ bl_0_29 br_0_29 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c29
*+ bl_0_29 br_0_29 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c29
+ bl_0_29 br_0_29 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c30
+ bl_0_30 br_0_30 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c30
*+ bl_0_30 br_0_30 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c30
*+ bl_0_30 br_0_30 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c30
*+ bl_0_30 br_0_30 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c30
*+ bl_0_30 br_0_30 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c30
*+ bl_0_30 br_0_30 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c30
*+ bl_0_30 br_0_30 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c30
*+ bl_0_30 br_0_30 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c30
*+ bl_0_30 br_0_30 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c30
*+ bl_0_30 br_0_30 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c30
*+ bl_0_30 br_0_30 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c30
*+ bl_0_30 br_0_30 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c30
*+ bl_0_30 br_0_30 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c30
*+ bl_0_30 br_0_30 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c30
*+ bl_0_30 br_0_30 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c30
*+ bl_0_30 br_0_30 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c30
*+ bl_0_30 br_0_30 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c30
*+ bl_0_30 br_0_30 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c30
*+ bl_0_30 br_0_30 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c30
*+ bl_0_30 br_0_30 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c30
*+ bl_0_30 br_0_30 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c30
*+ bl_0_30 br_0_30 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c30
*+ bl_0_30 br_0_30 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c30
*+ bl_0_30 br_0_30 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c30
*+ bl_0_30 br_0_30 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c30
*+ bl_0_30 br_0_30 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c30
*+ bl_0_30 br_0_30 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c30
*+ bl_0_30 br_0_30 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c30
*+ bl_0_30 br_0_30 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c30
*+ bl_0_30 br_0_30 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c30
*+ bl_0_30 br_0_30 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c30
*+ bl_0_30 br_0_30 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c30
*+ bl_0_30 br_0_30 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c30
*+ bl_0_30 br_0_30 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c30
*+ bl_0_30 br_0_30 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c30
*+ bl_0_30 br_0_30 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c30
*+ bl_0_30 br_0_30 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c30
*+ bl_0_30 br_0_30 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c30
*+ bl_0_30 br_0_30 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c30
*+ bl_0_30 br_0_30 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c30
*+ bl_0_30 br_0_30 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c30
*+ bl_0_30 br_0_30 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c30
*+ bl_0_30 br_0_30 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c30
*+ bl_0_30 br_0_30 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c30
*+ bl_0_30 br_0_30 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c30
*+ bl_0_30 br_0_30 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c30
*+ bl_0_30 br_0_30 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c30
*+ bl_0_30 br_0_30 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c30
*+ bl_0_30 br_0_30 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c30
*+ bl_0_30 br_0_30 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c30
*+ bl_0_30 br_0_30 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c30
*+ bl_0_30 br_0_30 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c30
*+ bl_0_30 br_0_30 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c30
*+ bl_0_30 br_0_30 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c30
*+ bl_0_30 br_0_30 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c30
*+ bl_0_30 br_0_30 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c30
*+ bl_0_30 br_0_30 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c30
*+ bl_0_30 br_0_30 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c30
*+ bl_0_30 br_0_30 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c30
*+ bl_0_30 br_0_30 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c30
*+ bl_0_30 br_0_30 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c30
*+ bl_0_30 br_0_30 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c30
*+ bl_0_30 br_0_30 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c30
*+ bl_0_30 br_0_30 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c30
*+ bl_0_30 br_0_30 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c30
*+ bl_0_30 br_0_30 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c30
*+ bl_0_30 br_0_30 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c30
*+ bl_0_30 br_0_30 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c30
*+ bl_0_30 br_0_30 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c30
*+ bl_0_30 br_0_30 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c30
*+ bl_0_30 br_0_30 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c30
*+ bl_0_30 br_0_30 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c30
*+ bl_0_30 br_0_30 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c30
*+ bl_0_30 br_0_30 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c30
*+ bl_0_30 br_0_30 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c30
*+ bl_0_30 br_0_30 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c30
*+ bl_0_30 br_0_30 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c30
*+ bl_0_30 br_0_30 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c30
*+ bl_0_30 br_0_30 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c30
*+ bl_0_30 br_0_30 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c30
*+ bl_0_30 br_0_30 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c30
*+ bl_0_30 br_0_30 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c30
*+ bl_0_30 br_0_30 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c30
*+ bl_0_30 br_0_30 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c30
*+ bl_0_30 br_0_30 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c30
*+ bl_0_30 br_0_30 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c30
*+ bl_0_30 br_0_30 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c30
*+ bl_0_30 br_0_30 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c30
*+ bl_0_30 br_0_30 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c30
*+ bl_0_30 br_0_30 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c30
*+ bl_0_30 br_0_30 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c30
*+ bl_0_30 br_0_30 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c30
*+ bl_0_30 br_0_30 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c30
*+ bl_0_30 br_0_30 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c30
*+ bl_0_30 br_0_30 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c30
*+ bl_0_30 br_0_30 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c30
*+ bl_0_30 br_0_30 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c30
*+ bl_0_30 br_0_30 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c30
*+ bl_0_30 br_0_30 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c30
*+ bl_0_30 br_0_30 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c30
*+ bl_0_30 br_0_30 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c30
*+ bl_0_30 br_0_30 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c30
*+ bl_0_30 br_0_30 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c30
*+ bl_0_30 br_0_30 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c30
*+ bl_0_30 br_0_30 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c30
*+ bl_0_30 br_0_30 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c30
*+ bl_0_30 br_0_30 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c30
*+ bl_0_30 br_0_30 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c30
*+ bl_0_30 br_0_30 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c30
*+ bl_0_30 br_0_30 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c30
*+ bl_0_30 br_0_30 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c30
*+ bl_0_30 br_0_30 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c30
*+ bl_0_30 br_0_30 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c30
*+ bl_0_30 br_0_30 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c30
*+ bl_0_30 br_0_30 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c30
*+ bl_0_30 br_0_30 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c30
*+ bl_0_30 br_0_30 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c30
*+ bl_0_30 br_0_30 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c30
*+ bl_0_30 br_0_30 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c30
*+ bl_0_30 br_0_30 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c30
*+ bl_0_30 br_0_30 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c30
*+ bl_0_30 br_0_30 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c30
*+ bl_0_30 br_0_30 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c30
*+ bl_0_30 br_0_30 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c30
*+ bl_0_30 br_0_30 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c30
*+ bl_0_30 br_0_30 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c30
*+ bl_0_30 br_0_30 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c30
+ bl_0_30 br_0_30 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c31
+ bl_0_31 br_0_31 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c31
*+ bl_0_31 br_0_31 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c31
*+ bl_0_31 br_0_31 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c31
*+ bl_0_31 br_0_31 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c31
*+ bl_0_31 br_0_31 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c31
*+ bl_0_31 br_0_31 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c31
*+ bl_0_31 br_0_31 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c31
*+ bl_0_31 br_0_31 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c31
*+ bl_0_31 br_0_31 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c31
*+ bl_0_31 br_0_31 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c31
*+ bl_0_31 br_0_31 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c31
*+ bl_0_31 br_0_31 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c31
*+ bl_0_31 br_0_31 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c31
*+ bl_0_31 br_0_31 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c31
*+ bl_0_31 br_0_31 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c31
*+ bl_0_31 br_0_31 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c31
*+ bl_0_31 br_0_31 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c31
*+ bl_0_31 br_0_31 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c31
*+ bl_0_31 br_0_31 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c31
*+ bl_0_31 br_0_31 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c31
*+ bl_0_31 br_0_31 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c31
*+ bl_0_31 br_0_31 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c31
*+ bl_0_31 br_0_31 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c31
*+ bl_0_31 br_0_31 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c31
*+ bl_0_31 br_0_31 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c31
*+ bl_0_31 br_0_31 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c31
*+ bl_0_31 br_0_31 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c31
*+ bl_0_31 br_0_31 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c31
*+ bl_0_31 br_0_31 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c31
*+ bl_0_31 br_0_31 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c31
*+ bl_0_31 br_0_31 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c31
*+ bl_0_31 br_0_31 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c31
*+ bl_0_31 br_0_31 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c31
*+ bl_0_31 br_0_31 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c31
*+ bl_0_31 br_0_31 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c31
*+ bl_0_31 br_0_31 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c31
*+ bl_0_31 br_0_31 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c31
*+ bl_0_31 br_0_31 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c31
*+ bl_0_31 br_0_31 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c31
*+ bl_0_31 br_0_31 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c31
*+ bl_0_31 br_0_31 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c31
*+ bl_0_31 br_0_31 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c31
*+ bl_0_31 br_0_31 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c31
*+ bl_0_31 br_0_31 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c31
*+ bl_0_31 br_0_31 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c31
*+ bl_0_31 br_0_31 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c31
*+ bl_0_31 br_0_31 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c31
*+ bl_0_31 br_0_31 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c31
*+ bl_0_31 br_0_31 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c31
*+ bl_0_31 br_0_31 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c31
*+ bl_0_31 br_0_31 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c31
*+ bl_0_31 br_0_31 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c31
*+ bl_0_31 br_0_31 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c31
*+ bl_0_31 br_0_31 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c31
*+ bl_0_31 br_0_31 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c31
*+ bl_0_31 br_0_31 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c31
*+ bl_0_31 br_0_31 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c31
*+ bl_0_31 br_0_31 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c31
*+ bl_0_31 br_0_31 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c31
*+ bl_0_31 br_0_31 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c31
*+ bl_0_31 br_0_31 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c31
*+ bl_0_31 br_0_31 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c31
*+ bl_0_31 br_0_31 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c31
*+ bl_0_31 br_0_31 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c31
*+ bl_0_31 br_0_31 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c31
*+ bl_0_31 br_0_31 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c31
*+ bl_0_31 br_0_31 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c31
*+ bl_0_31 br_0_31 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c31
*+ bl_0_31 br_0_31 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c31
*+ bl_0_31 br_0_31 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c31
*+ bl_0_31 br_0_31 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c31
*+ bl_0_31 br_0_31 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c31
*+ bl_0_31 br_0_31 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c31
*+ bl_0_31 br_0_31 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c31
*+ bl_0_31 br_0_31 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c31
*+ bl_0_31 br_0_31 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c31
*+ bl_0_31 br_0_31 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c31
*+ bl_0_31 br_0_31 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c31
*+ bl_0_31 br_0_31 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c31
*+ bl_0_31 br_0_31 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c31
*+ bl_0_31 br_0_31 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c31
*+ bl_0_31 br_0_31 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c31
*+ bl_0_31 br_0_31 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c31
*+ bl_0_31 br_0_31 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c31
*+ bl_0_31 br_0_31 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c31
*+ bl_0_31 br_0_31 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c31
*+ bl_0_31 br_0_31 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c31
*+ bl_0_31 br_0_31 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c31
*+ bl_0_31 br_0_31 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c31
*+ bl_0_31 br_0_31 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c31
*+ bl_0_31 br_0_31 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c31
*+ bl_0_31 br_0_31 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c31
*+ bl_0_31 br_0_31 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c31
*+ bl_0_31 br_0_31 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c31
*+ bl_0_31 br_0_31 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c31
*+ bl_0_31 br_0_31 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c31
*+ bl_0_31 br_0_31 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c31
*+ bl_0_31 br_0_31 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c31
*+ bl_0_31 br_0_31 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c31
*+ bl_0_31 br_0_31 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c31
*+ bl_0_31 br_0_31 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c31
*+ bl_0_31 br_0_31 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c31
*+ bl_0_31 br_0_31 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c31
*+ bl_0_31 br_0_31 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c31
*+ bl_0_31 br_0_31 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c31
*+ bl_0_31 br_0_31 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c31
*+ bl_0_31 br_0_31 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c31
*+ bl_0_31 br_0_31 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c31
*+ bl_0_31 br_0_31 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c31
*+ bl_0_31 br_0_31 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c31
*+ bl_0_31 br_0_31 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c31
*+ bl_0_31 br_0_31 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c31
*+ bl_0_31 br_0_31 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c31
*+ bl_0_31 br_0_31 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c31
*+ bl_0_31 br_0_31 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c31
*+ bl_0_31 br_0_31 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c31
*+ bl_0_31 br_0_31 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c31
*+ bl_0_31 br_0_31 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c31
*+ bl_0_31 br_0_31 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c31
*+ bl_0_31 br_0_31 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c31
*+ bl_0_31 br_0_31 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c31
*+ bl_0_31 br_0_31 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c31
*+ bl_0_31 br_0_31 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c31
*+ bl_0_31 br_0_31 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c31
*+ bl_0_31 br_0_31 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c31
*+ bl_0_31 br_0_31 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c31
*+ bl_0_31 br_0_31 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c31
+ bl_0_31 br_0_31 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c32
+ bl_0_32 br_0_32 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c32
*+ bl_0_32 br_0_32 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c32
*+ bl_0_32 br_0_32 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c32
*+ bl_0_32 br_0_32 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c32
*+ bl_0_32 br_0_32 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c32
*+ bl_0_32 br_0_32 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c32
*+ bl_0_32 br_0_32 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c32
*+ bl_0_32 br_0_32 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c32
*+ bl_0_32 br_0_32 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c32
*+ bl_0_32 br_0_32 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c32
*+ bl_0_32 br_0_32 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c32
*+ bl_0_32 br_0_32 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c32
*+ bl_0_32 br_0_32 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c32
*+ bl_0_32 br_0_32 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c32
*+ bl_0_32 br_0_32 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c32
*+ bl_0_32 br_0_32 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c32
*+ bl_0_32 br_0_32 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c32
*+ bl_0_32 br_0_32 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c32
*+ bl_0_32 br_0_32 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c32
*+ bl_0_32 br_0_32 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c32
*+ bl_0_32 br_0_32 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c32
*+ bl_0_32 br_0_32 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c32
*+ bl_0_32 br_0_32 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c32
*+ bl_0_32 br_0_32 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c32
*+ bl_0_32 br_0_32 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c32
*+ bl_0_32 br_0_32 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c32
*+ bl_0_32 br_0_32 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c32
*+ bl_0_32 br_0_32 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c32
*+ bl_0_32 br_0_32 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c32
*+ bl_0_32 br_0_32 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c32
*+ bl_0_32 br_0_32 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c32
*+ bl_0_32 br_0_32 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c32
*+ bl_0_32 br_0_32 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c32
*+ bl_0_32 br_0_32 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c32
*+ bl_0_32 br_0_32 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c32
*+ bl_0_32 br_0_32 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c32
*+ bl_0_32 br_0_32 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c32
*+ bl_0_32 br_0_32 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c32
*+ bl_0_32 br_0_32 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c32
*+ bl_0_32 br_0_32 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c32
*+ bl_0_32 br_0_32 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c32
*+ bl_0_32 br_0_32 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c32
*+ bl_0_32 br_0_32 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c32
*+ bl_0_32 br_0_32 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c32
*+ bl_0_32 br_0_32 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c32
*+ bl_0_32 br_0_32 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c32
*+ bl_0_32 br_0_32 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c32
*+ bl_0_32 br_0_32 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c32
*+ bl_0_32 br_0_32 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c32
*+ bl_0_32 br_0_32 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c32
*+ bl_0_32 br_0_32 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c32
*+ bl_0_32 br_0_32 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c32
*+ bl_0_32 br_0_32 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c32
*+ bl_0_32 br_0_32 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c32
*+ bl_0_32 br_0_32 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c32
*+ bl_0_32 br_0_32 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c32
*+ bl_0_32 br_0_32 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c32
*+ bl_0_32 br_0_32 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c32
*+ bl_0_32 br_0_32 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c32
*+ bl_0_32 br_0_32 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c32
*+ bl_0_32 br_0_32 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c32
*+ bl_0_32 br_0_32 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c32
*+ bl_0_32 br_0_32 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c32
*+ bl_0_32 br_0_32 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c32
*+ bl_0_32 br_0_32 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c32
*+ bl_0_32 br_0_32 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c32
*+ bl_0_32 br_0_32 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c32
*+ bl_0_32 br_0_32 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c32
*+ bl_0_32 br_0_32 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c32
*+ bl_0_32 br_0_32 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c32
*+ bl_0_32 br_0_32 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c32
*+ bl_0_32 br_0_32 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c32
*+ bl_0_32 br_0_32 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c32
*+ bl_0_32 br_0_32 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c32
*+ bl_0_32 br_0_32 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c32
*+ bl_0_32 br_0_32 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c32
*+ bl_0_32 br_0_32 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c32
*+ bl_0_32 br_0_32 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c32
*+ bl_0_32 br_0_32 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c32
*+ bl_0_32 br_0_32 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c32
*+ bl_0_32 br_0_32 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c32
*+ bl_0_32 br_0_32 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c32
*+ bl_0_32 br_0_32 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c32
*+ bl_0_32 br_0_32 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c32
*+ bl_0_32 br_0_32 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c32
*+ bl_0_32 br_0_32 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c32
*+ bl_0_32 br_0_32 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c32
*+ bl_0_32 br_0_32 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c32
*+ bl_0_32 br_0_32 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c32
*+ bl_0_32 br_0_32 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c32
*+ bl_0_32 br_0_32 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c32
*+ bl_0_32 br_0_32 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c32
*+ bl_0_32 br_0_32 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c32
*+ bl_0_32 br_0_32 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c32
*+ bl_0_32 br_0_32 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c32
*+ bl_0_32 br_0_32 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c32
*+ bl_0_32 br_0_32 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c32
*+ bl_0_32 br_0_32 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c32
*+ bl_0_32 br_0_32 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c32
*+ bl_0_32 br_0_32 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c32
*+ bl_0_32 br_0_32 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c32
*+ bl_0_32 br_0_32 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c32
*+ bl_0_32 br_0_32 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c32
*+ bl_0_32 br_0_32 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c32
*+ bl_0_32 br_0_32 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c32
*+ bl_0_32 br_0_32 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c32
*+ bl_0_32 br_0_32 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c32
*+ bl_0_32 br_0_32 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c32
*+ bl_0_32 br_0_32 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c32
*+ bl_0_32 br_0_32 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c32
*+ bl_0_32 br_0_32 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c32
*+ bl_0_32 br_0_32 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c32
*+ bl_0_32 br_0_32 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c32
*+ bl_0_32 br_0_32 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c32
*+ bl_0_32 br_0_32 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c32
*+ bl_0_32 br_0_32 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c32
*+ bl_0_32 br_0_32 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c32
*+ bl_0_32 br_0_32 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c32
*+ bl_0_32 br_0_32 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c32
*+ bl_0_32 br_0_32 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c32
*+ bl_0_32 br_0_32 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c32
*+ bl_0_32 br_0_32 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c32
*+ bl_0_32 br_0_32 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c32
*+ bl_0_32 br_0_32 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c32
*+ bl_0_32 br_0_32 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c32
*+ bl_0_32 br_0_32 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c32
*+ bl_0_32 br_0_32 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c32
+ bl_0_32 br_0_32 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c33
+ bl_0_33 br_0_33 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c33
*+ bl_0_33 br_0_33 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c33
*+ bl_0_33 br_0_33 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c33
*+ bl_0_33 br_0_33 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c33
*+ bl_0_33 br_0_33 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c33
*+ bl_0_33 br_0_33 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c33
*+ bl_0_33 br_0_33 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c33
*+ bl_0_33 br_0_33 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c33
*+ bl_0_33 br_0_33 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c33
*+ bl_0_33 br_0_33 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c33
*+ bl_0_33 br_0_33 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c33
*+ bl_0_33 br_0_33 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c33
*+ bl_0_33 br_0_33 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c33
*+ bl_0_33 br_0_33 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c33
*+ bl_0_33 br_0_33 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c33
*+ bl_0_33 br_0_33 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c33
*+ bl_0_33 br_0_33 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c33
*+ bl_0_33 br_0_33 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c33
*+ bl_0_33 br_0_33 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c33
*+ bl_0_33 br_0_33 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c33
*+ bl_0_33 br_0_33 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c33
*+ bl_0_33 br_0_33 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c33
*+ bl_0_33 br_0_33 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c33
*+ bl_0_33 br_0_33 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c33
*+ bl_0_33 br_0_33 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c33
*+ bl_0_33 br_0_33 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c33
*+ bl_0_33 br_0_33 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c33
*+ bl_0_33 br_0_33 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c33
*+ bl_0_33 br_0_33 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c33
*+ bl_0_33 br_0_33 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c33
*+ bl_0_33 br_0_33 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c33
*+ bl_0_33 br_0_33 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c33
*+ bl_0_33 br_0_33 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c33
*+ bl_0_33 br_0_33 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c33
*+ bl_0_33 br_0_33 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c33
*+ bl_0_33 br_0_33 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c33
*+ bl_0_33 br_0_33 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c33
*+ bl_0_33 br_0_33 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c33
*+ bl_0_33 br_0_33 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c33
*+ bl_0_33 br_0_33 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c33
*+ bl_0_33 br_0_33 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c33
*+ bl_0_33 br_0_33 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c33
*+ bl_0_33 br_0_33 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c33
*+ bl_0_33 br_0_33 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c33
*+ bl_0_33 br_0_33 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c33
*+ bl_0_33 br_0_33 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c33
*+ bl_0_33 br_0_33 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c33
*+ bl_0_33 br_0_33 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c33
*+ bl_0_33 br_0_33 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c33
*+ bl_0_33 br_0_33 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c33
*+ bl_0_33 br_0_33 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c33
*+ bl_0_33 br_0_33 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c33
*+ bl_0_33 br_0_33 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c33
*+ bl_0_33 br_0_33 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c33
*+ bl_0_33 br_0_33 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c33
*+ bl_0_33 br_0_33 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c33
*+ bl_0_33 br_0_33 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c33
*+ bl_0_33 br_0_33 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c33
*+ bl_0_33 br_0_33 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c33
*+ bl_0_33 br_0_33 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c33
*+ bl_0_33 br_0_33 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c33
*+ bl_0_33 br_0_33 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c33
*+ bl_0_33 br_0_33 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c33
*+ bl_0_33 br_0_33 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c33
*+ bl_0_33 br_0_33 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c33
*+ bl_0_33 br_0_33 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c33
*+ bl_0_33 br_0_33 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c33
*+ bl_0_33 br_0_33 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c33
*+ bl_0_33 br_0_33 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c33
*+ bl_0_33 br_0_33 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c33
*+ bl_0_33 br_0_33 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c33
*+ bl_0_33 br_0_33 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c33
*+ bl_0_33 br_0_33 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c33
*+ bl_0_33 br_0_33 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c33
*+ bl_0_33 br_0_33 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c33
*+ bl_0_33 br_0_33 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c33
*+ bl_0_33 br_0_33 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c33
*+ bl_0_33 br_0_33 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c33
*+ bl_0_33 br_0_33 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c33
*+ bl_0_33 br_0_33 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c33
*+ bl_0_33 br_0_33 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c33
*+ bl_0_33 br_0_33 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c33
*+ bl_0_33 br_0_33 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c33
*+ bl_0_33 br_0_33 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c33
*+ bl_0_33 br_0_33 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c33
*+ bl_0_33 br_0_33 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c33
*+ bl_0_33 br_0_33 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c33
*+ bl_0_33 br_0_33 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c33
*+ bl_0_33 br_0_33 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c33
*+ bl_0_33 br_0_33 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c33
*+ bl_0_33 br_0_33 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c33
*+ bl_0_33 br_0_33 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c33
*+ bl_0_33 br_0_33 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c33
*+ bl_0_33 br_0_33 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c33
*+ bl_0_33 br_0_33 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c33
*+ bl_0_33 br_0_33 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c33
*+ bl_0_33 br_0_33 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c33
*+ bl_0_33 br_0_33 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c33
*+ bl_0_33 br_0_33 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c33
*+ bl_0_33 br_0_33 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c33
*+ bl_0_33 br_0_33 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c33
*+ bl_0_33 br_0_33 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c33
*+ bl_0_33 br_0_33 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c33
*+ bl_0_33 br_0_33 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c33
*+ bl_0_33 br_0_33 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c33
*+ bl_0_33 br_0_33 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c33
*+ bl_0_33 br_0_33 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c33
*+ bl_0_33 br_0_33 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c33
*+ bl_0_33 br_0_33 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c33
*+ bl_0_33 br_0_33 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c33
*+ bl_0_33 br_0_33 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c33
*+ bl_0_33 br_0_33 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c33
*+ bl_0_33 br_0_33 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c33
*+ bl_0_33 br_0_33 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c33
*+ bl_0_33 br_0_33 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c33
*+ bl_0_33 br_0_33 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c33
*+ bl_0_33 br_0_33 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c33
*+ bl_0_33 br_0_33 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c33
*+ bl_0_33 br_0_33 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c33
*+ bl_0_33 br_0_33 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c33
*+ bl_0_33 br_0_33 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c33
*+ bl_0_33 br_0_33 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c33
*+ bl_0_33 br_0_33 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c33
*+ bl_0_33 br_0_33 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c33
*+ bl_0_33 br_0_33 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c33
*+ bl_0_33 br_0_33 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c33
*+ bl_0_33 br_0_33 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c33
+ bl_0_33 br_0_33 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c34
+ bl_0_34 br_0_34 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c34
*+ bl_0_34 br_0_34 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c34
*+ bl_0_34 br_0_34 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c34
*+ bl_0_34 br_0_34 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c34
*+ bl_0_34 br_0_34 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c34
*+ bl_0_34 br_0_34 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c34
*+ bl_0_34 br_0_34 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c34
*+ bl_0_34 br_0_34 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c34
*+ bl_0_34 br_0_34 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c34
*+ bl_0_34 br_0_34 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c34
*+ bl_0_34 br_0_34 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c34
*+ bl_0_34 br_0_34 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c34
*+ bl_0_34 br_0_34 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c34
*+ bl_0_34 br_0_34 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c34
*+ bl_0_34 br_0_34 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c34
*+ bl_0_34 br_0_34 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c34
*+ bl_0_34 br_0_34 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c34
*+ bl_0_34 br_0_34 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c34
*+ bl_0_34 br_0_34 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c34
*+ bl_0_34 br_0_34 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c34
*+ bl_0_34 br_0_34 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c34
*+ bl_0_34 br_0_34 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c34
*+ bl_0_34 br_0_34 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c34
*+ bl_0_34 br_0_34 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c34
*+ bl_0_34 br_0_34 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c34
*+ bl_0_34 br_0_34 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c34
*+ bl_0_34 br_0_34 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c34
*+ bl_0_34 br_0_34 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c34
*+ bl_0_34 br_0_34 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c34
*+ bl_0_34 br_0_34 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c34
*+ bl_0_34 br_0_34 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c34
*+ bl_0_34 br_0_34 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c34
*+ bl_0_34 br_0_34 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c34
*+ bl_0_34 br_0_34 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c34
*+ bl_0_34 br_0_34 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c34
*+ bl_0_34 br_0_34 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c34
*+ bl_0_34 br_0_34 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c34
*+ bl_0_34 br_0_34 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c34
*+ bl_0_34 br_0_34 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c34
*+ bl_0_34 br_0_34 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c34
*+ bl_0_34 br_0_34 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c34
*+ bl_0_34 br_0_34 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c34
*+ bl_0_34 br_0_34 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c34
*+ bl_0_34 br_0_34 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c34
*+ bl_0_34 br_0_34 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c34
*+ bl_0_34 br_0_34 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c34
*+ bl_0_34 br_0_34 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c34
*+ bl_0_34 br_0_34 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c34
*+ bl_0_34 br_0_34 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c34
*+ bl_0_34 br_0_34 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c34
*+ bl_0_34 br_0_34 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c34
*+ bl_0_34 br_0_34 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c34
*+ bl_0_34 br_0_34 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c34
*+ bl_0_34 br_0_34 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c34
*+ bl_0_34 br_0_34 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c34
*+ bl_0_34 br_0_34 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c34
*+ bl_0_34 br_0_34 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c34
*+ bl_0_34 br_0_34 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c34
*+ bl_0_34 br_0_34 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c34
*+ bl_0_34 br_0_34 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c34
*+ bl_0_34 br_0_34 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c34
*+ bl_0_34 br_0_34 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c34
*+ bl_0_34 br_0_34 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c34
*+ bl_0_34 br_0_34 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c34
*+ bl_0_34 br_0_34 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c34
*+ bl_0_34 br_0_34 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c34
*+ bl_0_34 br_0_34 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c34
*+ bl_0_34 br_0_34 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c34
*+ bl_0_34 br_0_34 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c34
*+ bl_0_34 br_0_34 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c34
*+ bl_0_34 br_0_34 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c34
*+ bl_0_34 br_0_34 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c34
*+ bl_0_34 br_0_34 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c34
*+ bl_0_34 br_0_34 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c34
*+ bl_0_34 br_0_34 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c34
*+ bl_0_34 br_0_34 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c34
*+ bl_0_34 br_0_34 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c34
*+ bl_0_34 br_0_34 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c34
*+ bl_0_34 br_0_34 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c34
*+ bl_0_34 br_0_34 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c34
*+ bl_0_34 br_0_34 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c34
*+ bl_0_34 br_0_34 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c34
*+ bl_0_34 br_0_34 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c34
*+ bl_0_34 br_0_34 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c34
*+ bl_0_34 br_0_34 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c34
*+ bl_0_34 br_0_34 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c34
*+ bl_0_34 br_0_34 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c34
*+ bl_0_34 br_0_34 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c34
*+ bl_0_34 br_0_34 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c34
*+ bl_0_34 br_0_34 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c34
*+ bl_0_34 br_0_34 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c34
*+ bl_0_34 br_0_34 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c34
*+ bl_0_34 br_0_34 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c34
*+ bl_0_34 br_0_34 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c34
*+ bl_0_34 br_0_34 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c34
*+ bl_0_34 br_0_34 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c34
*+ bl_0_34 br_0_34 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c34
*+ bl_0_34 br_0_34 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c34
*+ bl_0_34 br_0_34 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c34
*+ bl_0_34 br_0_34 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c34
*+ bl_0_34 br_0_34 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c34
*+ bl_0_34 br_0_34 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c34
*+ bl_0_34 br_0_34 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c34
*+ bl_0_34 br_0_34 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c34
*+ bl_0_34 br_0_34 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c34
*+ bl_0_34 br_0_34 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c34
*+ bl_0_34 br_0_34 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c34
*+ bl_0_34 br_0_34 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c34
*+ bl_0_34 br_0_34 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c34
*+ bl_0_34 br_0_34 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c34
*+ bl_0_34 br_0_34 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c34
*+ bl_0_34 br_0_34 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c34
*+ bl_0_34 br_0_34 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c34
*+ bl_0_34 br_0_34 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c34
*+ bl_0_34 br_0_34 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c34
*+ bl_0_34 br_0_34 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c34
*+ bl_0_34 br_0_34 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c34
*+ bl_0_34 br_0_34 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c34
*+ bl_0_34 br_0_34 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c34
*+ bl_0_34 br_0_34 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c34
*+ bl_0_34 br_0_34 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c34
*+ bl_0_34 br_0_34 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c34
*+ bl_0_34 br_0_34 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c34
*+ bl_0_34 br_0_34 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c34
*+ bl_0_34 br_0_34 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c34
*+ bl_0_34 br_0_34 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c34
*+ bl_0_34 br_0_34 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c34
+ bl_0_34 br_0_34 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c35
+ bl_0_35 br_0_35 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c35
*+ bl_0_35 br_0_35 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c35
*+ bl_0_35 br_0_35 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c35
*+ bl_0_35 br_0_35 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c35
*+ bl_0_35 br_0_35 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c35
*+ bl_0_35 br_0_35 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c35
*+ bl_0_35 br_0_35 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c35
*+ bl_0_35 br_0_35 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c35
*+ bl_0_35 br_0_35 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c35
*+ bl_0_35 br_0_35 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c35
*+ bl_0_35 br_0_35 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c35
*+ bl_0_35 br_0_35 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c35
*+ bl_0_35 br_0_35 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c35
*+ bl_0_35 br_0_35 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c35
*+ bl_0_35 br_0_35 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c35
*+ bl_0_35 br_0_35 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c35
*+ bl_0_35 br_0_35 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c35
*+ bl_0_35 br_0_35 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c35
*+ bl_0_35 br_0_35 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c35
*+ bl_0_35 br_0_35 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c35
*+ bl_0_35 br_0_35 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c35
*+ bl_0_35 br_0_35 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c35
*+ bl_0_35 br_0_35 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c35
*+ bl_0_35 br_0_35 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c35
*+ bl_0_35 br_0_35 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c35
*+ bl_0_35 br_0_35 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c35
*+ bl_0_35 br_0_35 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c35
*+ bl_0_35 br_0_35 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c35
*+ bl_0_35 br_0_35 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c35
*+ bl_0_35 br_0_35 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c35
*+ bl_0_35 br_0_35 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c35
*+ bl_0_35 br_0_35 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c35
*+ bl_0_35 br_0_35 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c35
*+ bl_0_35 br_0_35 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c35
*+ bl_0_35 br_0_35 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c35
*+ bl_0_35 br_0_35 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c35
*+ bl_0_35 br_0_35 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c35
*+ bl_0_35 br_0_35 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c35
*+ bl_0_35 br_0_35 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c35
*+ bl_0_35 br_0_35 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c35
*+ bl_0_35 br_0_35 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c35
*+ bl_0_35 br_0_35 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c35
*+ bl_0_35 br_0_35 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c35
*+ bl_0_35 br_0_35 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c35
*+ bl_0_35 br_0_35 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c35
*+ bl_0_35 br_0_35 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c35
*+ bl_0_35 br_0_35 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c35
*+ bl_0_35 br_0_35 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c35
*+ bl_0_35 br_0_35 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c35
*+ bl_0_35 br_0_35 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c35
*+ bl_0_35 br_0_35 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c35
*+ bl_0_35 br_0_35 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c35
*+ bl_0_35 br_0_35 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c35
*+ bl_0_35 br_0_35 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c35
*+ bl_0_35 br_0_35 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c35
*+ bl_0_35 br_0_35 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c35
*+ bl_0_35 br_0_35 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c35
*+ bl_0_35 br_0_35 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c35
*+ bl_0_35 br_0_35 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c35
*+ bl_0_35 br_0_35 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c35
*+ bl_0_35 br_0_35 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c35
*+ bl_0_35 br_0_35 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c35
*+ bl_0_35 br_0_35 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c35
*+ bl_0_35 br_0_35 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c35
*+ bl_0_35 br_0_35 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c35
*+ bl_0_35 br_0_35 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c35
*+ bl_0_35 br_0_35 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c35
*+ bl_0_35 br_0_35 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c35
*+ bl_0_35 br_0_35 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c35
*+ bl_0_35 br_0_35 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c35
*+ bl_0_35 br_0_35 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c35
*+ bl_0_35 br_0_35 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c35
*+ bl_0_35 br_0_35 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c35
*+ bl_0_35 br_0_35 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c35
*+ bl_0_35 br_0_35 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c35
*+ bl_0_35 br_0_35 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c35
*+ bl_0_35 br_0_35 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c35
*+ bl_0_35 br_0_35 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c35
*+ bl_0_35 br_0_35 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c35
*+ bl_0_35 br_0_35 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c35
*+ bl_0_35 br_0_35 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c35
*+ bl_0_35 br_0_35 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c35
*+ bl_0_35 br_0_35 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c35
*+ bl_0_35 br_0_35 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c35
*+ bl_0_35 br_0_35 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c35
*+ bl_0_35 br_0_35 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c35
*+ bl_0_35 br_0_35 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c35
*+ bl_0_35 br_0_35 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c35
*+ bl_0_35 br_0_35 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c35
*+ bl_0_35 br_0_35 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c35
*+ bl_0_35 br_0_35 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c35
*+ bl_0_35 br_0_35 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c35
*+ bl_0_35 br_0_35 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c35
*+ bl_0_35 br_0_35 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c35
*+ bl_0_35 br_0_35 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c35
*+ bl_0_35 br_0_35 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c35
*+ bl_0_35 br_0_35 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c35
*+ bl_0_35 br_0_35 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c35
*+ bl_0_35 br_0_35 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c35
*+ bl_0_35 br_0_35 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c35
*+ bl_0_35 br_0_35 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c35
*+ bl_0_35 br_0_35 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c35
*+ bl_0_35 br_0_35 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c35
*+ bl_0_35 br_0_35 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c35
*+ bl_0_35 br_0_35 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c35
*+ bl_0_35 br_0_35 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c35
*+ bl_0_35 br_0_35 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c35
*+ bl_0_35 br_0_35 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c35
*+ bl_0_35 br_0_35 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c35
*+ bl_0_35 br_0_35 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c35
*+ bl_0_35 br_0_35 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c35
*+ bl_0_35 br_0_35 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c35
*+ bl_0_35 br_0_35 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c35
*+ bl_0_35 br_0_35 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c35
*+ bl_0_35 br_0_35 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c35
*+ bl_0_35 br_0_35 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c35
*+ bl_0_35 br_0_35 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c35
*+ bl_0_35 br_0_35 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c35
*+ bl_0_35 br_0_35 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c35
*+ bl_0_35 br_0_35 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c35
*+ bl_0_35 br_0_35 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c35
*+ bl_0_35 br_0_35 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c35
*+ bl_0_35 br_0_35 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c35
*+ bl_0_35 br_0_35 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c35
*+ bl_0_35 br_0_35 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c35
*+ bl_0_35 br_0_35 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c35
*+ bl_0_35 br_0_35 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c35
+ bl_0_35 br_0_35 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c36
+ bl_0_36 br_0_36 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c36
*+ bl_0_36 br_0_36 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c36
*+ bl_0_36 br_0_36 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c36
*+ bl_0_36 br_0_36 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c36
*+ bl_0_36 br_0_36 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c36
*+ bl_0_36 br_0_36 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c36
*+ bl_0_36 br_0_36 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c36
*+ bl_0_36 br_0_36 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c36
*+ bl_0_36 br_0_36 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c36
*+ bl_0_36 br_0_36 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c36
*+ bl_0_36 br_0_36 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c36
*+ bl_0_36 br_0_36 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c36
*+ bl_0_36 br_0_36 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c36
*+ bl_0_36 br_0_36 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c36
*+ bl_0_36 br_0_36 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c36
*+ bl_0_36 br_0_36 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c36
*+ bl_0_36 br_0_36 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c36
*+ bl_0_36 br_0_36 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c36
*+ bl_0_36 br_0_36 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c36
*+ bl_0_36 br_0_36 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c36
*+ bl_0_36 br_0_36 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c36
*+ bl_0_36 br_0_36 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c36
*+ bl_0_36 br_0_36 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c36
*+ bl_0_36 br_0_36 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c36
*+ bl_0_36 br_0_36 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c36
*+ bl_0_36 br_0_36 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c36
*+ bl_0_36 br_0_36 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c36
*+ bl_0_36 br_0_36 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c36
*+ bl_0_36 br_0_36 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c36
*+ bl_0_36 br_0_36 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c36
*+ bl_0_36 br_0_36 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c36
*+ bl_0_36 br_0_36 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c36
*+ bl_0_36 br_0_36 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c36
*+ bl_0_36 br_0_36 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c36
*+ bl_0_36 br_0_36 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c36
*+ bl_0_36 br_0_36 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c36
*+ bl_0_36 br_0_36 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c36
*+ bl_0_36 br_0_36 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c36
*+ bl_0_36 br_0_36 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c36
*+ bl_0_36 br_0_36 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c36
*+ bl_0_36 br_0_36 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c36
*+ bl_0_36 br_0_36 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c36
*+ bl_0_36 br_0_36 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c36
*+ bl_0_36 br_0_36 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c36
*+ bl_0_36 br_0_36 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c36
*+ bl_0_36 br_0_36 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c36
*+ bl_0_36 br_0_36 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c36
*+ bl_0_36 br_0_36 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c36
*+ bl_0_36 br_0_36 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c36
*+ bl_0_36 br_0_36 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c36
*+ bl_0_36 br_0_36 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c36
*+ bl_0_36 br_0_36 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c36
*+ bl_0_36 br_0_36 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c36
*+ bl_0_36 br_0_36 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c36
*+ bl_0_36 br_0_36 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c36
*+ bl_0_36 br_0_36 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c36
*+ bl_0_36 br_0_36 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c36
*+ bl_0_36 br_0_36 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c36
*+ bl_0_36 br_0_36 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c36
*+ bl_0_36 br_0_36 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c36
*+ bl_0_36 br_0_36 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c36
*+ bl_0_36 br_0_36 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c36
*+ bl_0_36 br_0_36 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c36
*+ bl_0_36 br_0_36 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c36
*+ bl_0_36 br_0_36 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c36
*+ bl_0_36 br_0_36 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c36
*+ bl_0_36 br_0_36 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c36
*+ bl_0_36 br_0_36 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c36
*+ bl_0_36 br_0_36 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c36
*+ bl_0_36 br_0_36 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c36
*+ bl_0_36 br_0_36 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c36
*+ bl_0_36 br_0_36 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c36
*+ bl_0_36 br_0_36 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c36
*+ bl_0_36 br_0_36 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c36
*+ bl_0_36 br_0_36 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c36
*+ bl_0_36 br_0_36 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c36
*+ bl_0_36 br_0_36 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c36
*+ bl_0_36 br_0_36 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c36
*+ bl_0_36 br_0_36 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c36
*+ bl_0_36 br_0_36 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c36
*+ bl_0_36 br_0_36 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c36
*+ bl_0_36 br_0_36 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c36
*+ bl_0_36 br_0_36 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c36
*+ bl_0_36 br_0_36 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c36
*+ bl_0_36 br_0_36 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c36
*+ bl_0_36 br_0_36 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c36
*+ bl_0_36 br_0_36 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c36
*+ bl_0_36 br_0_36 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c36
*+ bl_0_36 br_0_36 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c36
*+ bl_0_36 br_0_36 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c36
*+ bl_0_36 br_0_36 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c36
*+ bl_0_36 br_0_36 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c36
*+ bl_0_36 br_0_36 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c36
*+ bl_0_36 br_0_36 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c36
*+ bl_0_36 br_0_36 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c36
*+ bl_0_36 br_0_36 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c36
*+ bl_0_36 br_0_36 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c36
*+ bl_0_36 br_0_36 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c36
*+ bl_0_36 br_0_36 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c36
*+ bl_0_36 br_0_36 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c36
*+ bl_0_36 br_0_36 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c36
*+ bl_0_36 br_0_36 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c36
*+ bl_0_36 br_0_36 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c36
*+ bl_0_36 br_0_36 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c36
*+ bl_0_36 br_0_36 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c36
*+ bl_0_36 br_0_36 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c36
*+ bl_0_36 br_0_36 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c36
*+ bl_0_36 br_0_36 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c36
*+ bl_0_36 br_0_36 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c36
*+ bl_0_36 br_0_36 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c36
*+ bl_0_36 br_0_36 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c36
*+ bl_0_36 br_0_36 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c36
*+ bl_0_36 br_0_36 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c36
*+ bl_0_36 br_0_36 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c36
*+ bl_0_36 br_0_36 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c36
*+ bl_0_36 br_0_36 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c36
*+ bl_0_36 br_0_36 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c36
*+ bl_0_36 br_0_36 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c36
*+ bl_0_36 br_0_36 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c36
*+ bl_0_36 br_0_36 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c36
*+ bl_0_36 br_0_36 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c36
*+ bl_0_36 br_0_36 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c36
*+ bl_0_36 br_0_36 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c36
*+ bl_0_36 br_0_36 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c36
*+ bl_0_36 br_0_36 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c36
*+ bl_0_36 br_0_36 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c36
*+ bl_0_36 br_0_36 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c36
+ bl_0_36 br_0_36 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c37
+ bl_0_37 br_0_37 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c37
*+ bl_0_37 br_0_37 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c37
*+ bl_0_37 br_0_37 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c37
*+ bl_0_37 br_0_37 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c37
*+ bl_0_37 br_0_37 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c37
*+ bl_0_37 br_0_37 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c37
*+ bl_0_37 br_0_37 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c37
*+ bl_0_37 br_0_37 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c37
*+ bl_0_37 br_0_37 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c37
*+ bl_0_37 br_0_37 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c37
*+ bl_0_37 br_0_37 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c37
*+ bl_0_37 br_0_37 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c37
*+ bl_0_37 br_0_37 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c37
*+ bl_0_37 br_0_37 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c37
*+ bl_0_37 br_0_37 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c37
*+ bl_0_37 br_0_37 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c37
*+ bl_0_37 br_0_37 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c37
*+ bl_0_37 br_0_37 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c37
*+ bl_0_37 br_0_37 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c37
*+ bl_0_37 br_0_37 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c37
*+ bl_0_37 br_0_37 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c37
*+ bl_0_37 br_0_37 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c37
*+ bl_0_37 br_0_37 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c37
*+ bl_0_37 br_0_37 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c37
*+ bl_0_37 br_0_37 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c37
*+ bl_0_37 br_0_37 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c37
*+ bl_0_37 br_0_37 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c37
*+ bl_0_37 br_0_37 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c37
*+ bl_0_37 br_0_37 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c37
*+ bl_0_37 br_0_37 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c37
*+ bl_0_37 br_0_37 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c37
*+ bl_0_37 br_0_37 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c37
*+ bl_0_37 br_0_37 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c37
*+ bl_0_37 br_0_37 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c37
*+ bl_0_37 br_0_37 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c37
*+ bl_0_37 br_0_37 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c37
*+ bl_0_37 br_0_37 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c37
*+ bl_0_37 br_0_37 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c37
*+ bl_0_37 br_0_37 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c37
*+ bl_0_37 br_0_37 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c37
*+ bl_0_37 br_0_37 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c37
*+ bl_0_37 br_0_37 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c37
*+ bl_0_37 br_0_37 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c37
*+ bl_0_37 br_0_37 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c37
*+ bl_0_37 br_0_37 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c37
*+ bl_0_37 br_0_37 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c37
*+ bl_0_37 br_0_37 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c37
*+ bl_0_37 br_0_37 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c37
*+ bl_0_37 br_0_37 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c37
*+ bl_0_37 br_0_37 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c37
*+ bl_0_37 br_0_37 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c37
*+ bl_0_37 br_0_37 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c37
*+ bl_0_37 br_0_37 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c37
*+ bl_0_37 br_0_37 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c37
*+ bl_0_37 br_0_37 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c37
*+ bl_0_37 br_0_37 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c37
*+ bl_0_37 br_0_37 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c37
*+ bl_0_37 br_0_37 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c37
*+ bl_0_37 br_0_37 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c37
*+ bl_0_37 br_0_37 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c37
*+ bl_0_37 br_0_37 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c37
*+ bl_0_37 br_0_37 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c37
*+ bl_0_37 br_0_37 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c37
*+ bl_0_37 br_0_37 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c37
*+ bl_0_37 br_0_37 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c37
*+ bl_0_37 br_0_37 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c37
*+ bl_0_37 br_0_37 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c37
*+ bl_0_37 br_0_37 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c37
*+ bl_0_37 br_0_37 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c37
*+ bl_0_37 br_0_37 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c37
*+ bl_0_37 br_0_37 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c37
*+ bl_0_37 br_0_37 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c37
*+ bl_0_37 br_0_37 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c37
*+ bl_0_37 br_0_37 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c37
*+ bl_0_37 br_0_37 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c37
*+ bl_0_37 br_0_37 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c37
*+ bl_0_37 br_0_37 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c37
*+ bl_0_37 br_0_37 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c37
*+ bl_0_37 br_0_37 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c37
*+ bl_0_37 br_0_37 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c37
*+ bl_0_37 br_0_37 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c37
*+ bl_0_37 br_0_37 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c37
*+ bl_0_37 br_0_37 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c37
*+ bl_0_37 br_0_37 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c37
*+ bl_0_37 br_0_37 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c37
*+ bl_0_37 br_0_37 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c37
*+ bl_0_37 br_0_37 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c37
*+ bl_0_37 br_0_37 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c37
*+ bl_0_37 br_0_37 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c37
*+ bl_0_37 br_0_37 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c37
*+ bl_0_37 br_0_37 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c37
*+ bl_0_37 br_0_37 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c37
*+ bl_0_37 br_0_37 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c37
*+ bl_0_37 br_0_37 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c37
*+ bl_0_37 br_0_37 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c37
*+ bl_0_37 br_0_37 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c37
*+ bl_0_37 br_0_37 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c37
*+ bl_0_37 br_0_37 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c37
*+ bl_0_37 br_0_37 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c37
*+ bl_0_37 br_0_37 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c37
*+ bl_0_37 br_0_37 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c37
*+ bl_0_37 br_0_37 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c37
*+ bl_0_37 br_0_37 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c37
*+ bl_0_37 br_0_37 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c37
*+ bl_0_37 br_0_37 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c37
*+ bl_0_37 br_0_37 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c37
*+ bl_0_37 br_0_37 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c37
*+ bl_0_37 br_0_37 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c37
*+ bl_0_37 br_0_37 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c37
*+ bl_0_37 br_0_37 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c37
*+ bl_0_37 br_0_37 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c37
*+ bl_0_37 br_0_37 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c37
*+ bl_0_37 br_0_37 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c37
*+ bl_0_37 br_0_37 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c37
*+ bl_0_37 br_0_37 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c37
*+ bl_0_37 br_0_37 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c37
*+ bl_0_37 br_0_37 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c37
*+ bl_0_37 br_0_37 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c37
*+ bl_0_37 br_0_37 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c37
*+ bl_0_37 br_0_37 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c37
*+ bl_0_37 br_0_37 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c37
*+ bl_0_37 br_0_37 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c37
*+ bl_0_37 br_0_37 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c37
*+ bl_0_37 br_0_37 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c37
*+ bl_0_37 br_0_37 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c37
*+ bl_0_37 br_0_37 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c37
*+ bl_0_37 br_0_37 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c37
+ bl_0_37 br_0_37 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c38
+ bl_0_38 br_0_38 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c38
*+ bl_0_38 br_0_38 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c38
*+ bl_0_38 br_0_38 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c38
*+ bl_0_38 br_0_38 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c38
*+ bl_0_38 br_0_38 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c38
*+ bl_0_38 br_0_38 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c38
*+ bl_0_38 br_0_38 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c38
*+ bl_0_38 br_0_38 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c38
*+ bl_0_38 br_0_38 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c38
*+ bl_0_38 br_0_38 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c38
*+ bl_0_38 br_0_38 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c38
*+ bl_0_38 br_0_38 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c38
*+ bl_0_38 br_0_38 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c38
*+ bl_0_38 br_0_38 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c38
*+ bl_0_38 br_0_38 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c38
*+ bl_0_38 br_0_38 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c38
*+ bl_0_38 br_0_38 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c38
*+ bl_0_38 br_0_38 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c38
*+ bl_0_38 br_0_38 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c38
*+ bl_0_38 br_0_38 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c38
*+ bl_0_38 br_0_38 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c38
*+ bl_0_38 br_0_38 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c38
*+ bl_0_38 br_0_38 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c38
*+ bl_0_38 br_0_38 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c38
*+ bl_0_38 br_0_38 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c38
*+ bl_0_38 br_0_38 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c38
*+ bl_0_38 br_0_38 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c38
*+ bl_0_38 br_0_38 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c38
*+ bl_0_38 br_0_38 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c38
*+ bl_0_38 br_0_38 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c38
*+ bl_0_38 br_0_38 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c38
*+ bl_0_38 br_0_38 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c38
*+ bl_0_38 br_0_38 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c38
*+ bl_0_38 br_0_38 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c38
*+ bl_0_38 br_0_38 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c38
*+ bl_0_38 br_0_38 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c38
*+ bl_0_38 br_0_38 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c38
*+ bl_0_38 br_0_38 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c38
*+ bl_0_38 br_0_38 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c38
*+ bl_0_38 br_0_38 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c38
*+ bl_0_38 br_0_38 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c38
*+ bl_0_38 br_0_38 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c38
*+ bl_0_38 br_0_38 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c38
*+ bl_0_38 br_0_38 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c38
*+ bl_0_38 br_0_38 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c38
*+ bl_0_38 br_0_38 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c38
*+ bl_0_38 br_0_38 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c38
*+ bl_0_38 br_0_38 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c38
*+ bl_0_38 br_0_38 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c38
*+ bl_0_38 br_0_38 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c38
*+ bl_0_38 br_0_38 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c38
*+ bl_0_38 br_0_38 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c38
*+ bl_0_38 br_0_38 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c38
*+ bl_0_38 br_0_38 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c38
*+ bl_0_38 br_0_38 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c38
*+ bl_0_38 br_0_38 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c38
*+ bl_0_38 br_0_38 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c38
*+ bl_0_38 br_0_38 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c38
*+ bl_0_38 br_0_38 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c38
*+ bl_0_38 br_0_38 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c38
*+ bl_0_38 br_0_38 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c38
*+ bl_0_38 br_0_38 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c38
*+ bl_0_38 br_0_38 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c38
*+ bl_0_38 br_0_38 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c38
*+ bl_0_38 br_0_38 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c38
*+ bl_0_38 br_0_38 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c38
*+ bl_0_38 br_0_38 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c38
*+ bl_0_38 br_0_38 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c38
*+ bl_0_38 br_0_38 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c38
*+ bl_0_38 br_0_38 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c38
*+ bl_0_38 br_0_38 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c38
*+ bl_0_38 br_0_38 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c38
*+ bl_0_38 br_0_38 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c38
*+ bl_0_38 br_0_38 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c38
*+ bl_0_38 br_0_38 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c38
*+ bl_0_38 br_0_38 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c38
*+ bl_0_38 br_0_38 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c38
*+ bl_0_38 br_0_38 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c38
*+ bl_0_38 br_0_38 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c38
*+ bl_0_38 br_0_38 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c38
*+ bl_0_38 br_0_38 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c38
*+ bl_0_38 br_0_38 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c38
*+ bl_0_38 br_0_38 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c38
*+ bl_0_38 br_0_38 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c38
*+ bl_0_38 br_0_38 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c38
*+ bl_0_38 br_0_38 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c38
*+ bl_0_38 br_0_38 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c38
*+ bl_0_38 br_0_38 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c38
*+ bl_0_38 br_0_38 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c38
*+ bl_0_38 br_0_38 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c38
*+ bl_0_38 br_0_38 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c38
*+ bl_0_38 br_0_38 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c38
*+ bl_0_38 br_0_38 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c38
*+ bl_0_38 br_0_38 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c38
*+ bl_0_38 br_0_38 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c38
*+ bl_0_38 br_0_38 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c38
*+ bl_0_38 br_0_38 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c38
*+ bl_0_38 br_0_38 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c38
*+ bl_0_38 br_0_38 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c38
*+ bl_0_38 br_0_38 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c38
*+ bl_0_38 br_0_38 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c38
*+ bl_0_38 br_0_38 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c38
*+ bl_0_38 br_0_38 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c38
*+ bl_0_38 br_0_38 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c38
*+ bl_0_38 br_0_38 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c38
*+ bl_0_38 br_0_38 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c38
*+ bl_0_38 br_0_38 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c38
*+ bl_0_38 br_0_38 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c38
*+ bl_0_38 br_0_38 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c38
*+ bl_0_38 br_0_38 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c38
*+ bl_0_38 br_0_38 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c38
*+ bl_0_38 br_0_38 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c38
*+ bl_0_38 br_0_38 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c38
*+ bl_0_38 br_0_38 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c38
*+ bl_0_38 br_0_38 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c38
*+ bl_0_38 br_0_38 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c38
*+ bl_0_38 br_0_38 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c38
*+ bl_0_38 br_0_38 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c38
*+ bl_0_38 br_0_38 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c38
*+ bl_0_38 br_0_38 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c38
*+ bl_0_38 br_0_38 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c38
*+ bl_0_38 br_0_38 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c38
*+ bl_0_38 br_0_38 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c38
*+ bl_0_38 br_0_38 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c38
*+ bl_0_38 br_0_38 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c38
*+ bl_0_38 br_0_38 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c38
*+ bl_0_38 br_0_38 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c38
+ bl_0_38 br_0_38 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c39
+ bl_0_39 br_0_39 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c39
*+ bl_0_39 br_0_39 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c39
*+ bl_0_39 br_0_39 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c39
*+ bl_0_39 br_0_39 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c39
*+ bl_0_39 br_0_39 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c39
*+ bl_0_39 br_0_39 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c39
*+ bl_0_39 br_0_39 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c39
*+ bl_0_39 br_0_39 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c39
*+ bl_0_39 br_0_39 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c39
*+ bl_0_39 br_0_39 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c39
*+ bl_0_39 br_0_39 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c39
*+ bl_0_39 br_0_39 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c39
*+ bl_0_39 br_0_39 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c39
*+ bl_0_39 br_0_39 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c39
*+ bl_0_39 br_0_39 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c39
*+ bl_0_39 br_0_39 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c39
*+ bl_0_39 br_0_39 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c39
*+ bl_0_39 br_0_39 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c39
*+ bl_0_39 br_0_39 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c39
*+ bl_0_39 br_0_39 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c39
*+ bl_0_39 br_0_39 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c39
*+ bl_0_39 br_0_39 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c39
*+ bl_0_39 br_0_39 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c39
*+ bl_0_39 br_0_39 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c39
*+ bl_0_39 br_0_39 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c39
*+ bl_0_39 br_0_39 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c39
*+ bl_0_39 br_0_39 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c39
*+ bl_0_39 br_0_39 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c39
*+ bl_0_39 br_0_39 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c39
*+ bl_0_39 br_0_39 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c39
*+ bl_0_39 br_0_39 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c39
*+ bl_0_39 br_0_39 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c39
*+ bl_0_39 br_0_39 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c39
*+ bl_0_39 br_0_39 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c39
*+ bl_0_39 br_0_39 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c39
*+ bl_0_39 br_0_39 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c39
*+ bl_0_39 br_0_39 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c39
*+ bl_0_39 br_0_39 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c39
*+ bl_0_39 br_0_39 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c39
*+ bl_0_39 br_0_39 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c39
*+ bl_0_39 br_0_39 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c39
*+ bl_0_39 br_0_39 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c39
*+ bl_0_39 br_0_39 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c39
*+ bl_0_39 br_0_39 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c39
*+ bl_0_39 br_0_39 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c39
*+ bl_0_39 br_0_39 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c39
*+ bl_0_39 br_0_39 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c39
*+ bl_0_39 br_0_39 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c39
*+ bl_0_39 br_0_39 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c39
*+ bl_0_39 br_0_39 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c39
*+ bl_0_39 br_0_39 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c39
*+ bl_0_39 br_0_39 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c39
*+ bl_0_39 br_0_39 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c39
*+ bl_0_39 br_0_39 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c39
*+ bl_0_39 br_0_39 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c39
*+ bl_0_39 br_0_39 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c39
*+ bl_0_39 br_0_39 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c39
*+ bl_0_39 br_0_39 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c39
*+ bl_0_39 br_0_39 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c39
*+ bl_0_39 br_0_39 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c39
*+ bl_0_39 br_0_39 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c39
*+ bl_0_39 br_0_39 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c39
*+ bl_0_39 br_0_39 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c39
*+ bl_0_39 br_0_39 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c39
*+ bl_0_39 br_0_39 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c39
*+ bl_0_39 br_0_39 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c39
*+ bl_0_39 br_0_39 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c39
*+ bl_0_39 br_0_39 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c39
*+ bl_0_39 br_0_39 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c39
*+ bl_0_39 br_0_39 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c39
*+ bl_0_39 br_0_39 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c39
*+ bl_0_39 br_0_39 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c39
*+ bl_0_39 br_0_39 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c39
*+ bl_0_39 br_0_39 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c39
*+ bl_0_39 br_0_39 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c39
*+ bl_0_39 br_0_39 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c39
*+ bl_0_39 br_0_39 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c39
*+ bl_0_39 br_0_39 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c39
*+ bl_0_39 br_0_39 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c39
*+ bl_0_39 br_0_39 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c39
*+ bl_0_39 br_0_39 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c39
*+ bl_0_39 br_0_39 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c39
*+ bl_0_39 br_0_39 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c39
*+ bl_0_39 br_0_39 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c39
*+ bl_0_39 br_0_39 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c39
*+ bl_0_39 br_0_39 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c39
*+ bl_0_39 br_0_39 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c39
*+ bl_0_39 br_0_39 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c39
*+ bl_0_39 br_0_39 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c39
*+ bl_0_39 br_0_39 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c39
*+ bl_0_39 br_0_39 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c39
*+ bl_0_39 br_0_39 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c39
*+ bl_0_39 br_0_39 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c39
*+ bl_0_39 br_0_39 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c39
*+ bl_0_39 br_0_39 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c39
*+ bl_0_39 br_0_39 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c39
*+ bl_0_39 br_0_39 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c39
*+ bl_0_39 br_0_39 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c39
*+ bl_0_39 br_0_39 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c39
*+ bl_0_39 br_0_39 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c39
*+ bl_0_39 br_0_39 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c39
*+ bl_0_39 br_0_39 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c39
*+ bl_0_39 br_0_39 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c39
*+ bl_0_39 br_0_39 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c39
*+ bl_0_39 br_0_39 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c39
*+ bl_0_39 br_0_39 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c39
*+ bl_0_39 br_0_39 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c39
*+ bl_0_39 br_0_39 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c39
*+ bl_0_39 br_0_39 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c39
*+ bl_0_39 br_0_39 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c39
*+ bl_0_39 br_0_39 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c39
*+ bl_0_39 br_0_39 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c39
*+ bl_0_39 br_0_39 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c39
*+ bl_0_39 br_0_39 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c39
*+ bl_0_39 br_0_39 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c39
*+ bl_0_39 br_0_39 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c39
*+ bl_0_39 br_0_39 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c39
*+ bl_0_39 br_0_39 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c39
*+ bl_0_39 br_0_39 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c39
*+ bl_0_39 br_0_39 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c39
*+ bl_0_39 br_0_39 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c39
*+ bl_0_39 br_0_39 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c39
*+ bl_0_39 br_0_39 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c39
*+ bl_0_39 br_0_39 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c39
*+ bl_0_39 br_0_39 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c39
*+ bl_0_39 br_0_39 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c39
*+ bl_0_39 br_0_39 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c39
+ bl_0_39 br_0_39 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c40
+ bl_0_40 br_0_40 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c40
*+ bl_0_40 br_0_40 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c40
*+ bl_0_40 br_0_40 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c40
*+ bl_0_40 br_0_40 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c40
*+ bl_0_40 br_0_40 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c40
*+ bl_0_40 br_0_40 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c40
*+ bl_0_40 br_0_40 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c40
*+ bl_0_40 br_0_40 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c40
*+ bl_0_40 br_0_40 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c40
*+ bl_0_40 br_0_40 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c40
*+ bl_0_40 br_0_40 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c40
*+ bl_0_40 br_0_40 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c40
*+ bl_0_40 br_0_40 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c40
*+ bl_0_40 br_0_40 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c40
*+ bl_0_40 br_0_40 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c40
*+ bl_0_40 br_0_40 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c40
*+ bl_0_40 br_0_40 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c40
*+ bl_0_40 br_0_40 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c40
*+ bl_0_40 br_0_40 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c40
*+ bl_0_40 br_0_40 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c40
*+ bl_0_40 br_0_40 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c40
*+ bl_0_40 br_0_40 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c40
*+ bl_0_40 br_0_40 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c40
*+ bl_0_40 br_0_40 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c40
*+ bl_0_40 br_0_40 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c40
*+ bl_0_40 br_0_40 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c40
*+ bl_0_40 br_0_40 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c40
*+ bl_0_40 br_0_40 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c40
*+ bl_0_40 br_0_40 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c40
*+ bl_0_40 br_0_40 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c40
*+ bl_0_40 br_0_40 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c40
*+ bl_0_40 br_0_40 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c40
*+ bl_0_40 br_0_40 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c40
*+ bl_0_40 br_0_40 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c40
*+ bl_0_40 br_0_40 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c40
*+ bl_0_40 br_0_40 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c40
*+ bl_0_40 br_0_40 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c40
*+ bl_0_40 br_0_40 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c40
*+ bl_0_40 br_0_40 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c40
*+ bl_0_40 br_0_40 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c40
*+ bl_0_40 br_0_40 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c40
*+ bl_0_40 br_0_40 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c40
*+ bl_0_40 br_0_40 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c40
*+ bl_0_40 br_0_40 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c40
*+ bl_0_40 br_0_40 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c40
*+ bl_0_40 br_0_40 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c40
*+ bl_0_40 br_0_40 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c40
*+ bl_0_40 br_0_40 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c40
*+ bl_0_40 br_0_40 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c40
*+ bl_0_40 br_0_40 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c40
*+ bl_0_40 br_0_40 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c40
*+ bl_0_40 br_0_40 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c40
*+ bl_0_40 br_0_40 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c40
*+ bl_0_40 br_0_40 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c40
*+ bl_0_40 br_0_40 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c40
*+ bl_0_40 br_0_40 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c40
*+ bl_0_40 br_0_40 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c40
*+ bl_0_40 br_0_40 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c40
*+ bl_0_40 br_0_40 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c40
*+ bl_0_40 br_0_40 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c40
*+ bl_0_40 br_0_40 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c40
*+ bl_0_40 br_0_40 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c40
*+ bl_0_40 br_0_40 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c40
*+ bl_0_40 br_0_40 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c40
*+ bl_0_40 br_0_40 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c40
*+ bl_0_40 br_0_40 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c40
*+ bl_0_40 br_0_40 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c40
*+ bl_0_40 br_0_40 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c40
*+ bl_0_40 br_0_40 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c40
*+ bl_0_40 br_0_40 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c40
*+ bl_0_40 br_0_40 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c40
*+ bl_0_40 br_0_40 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c40
*+ bl_0_40 br_0_40 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c40
*+ bl_0_40 br_0_40 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c40
*+ bl_0_40 br_0_40 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c40
*+ bl_0_40 br_0_40 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c40
*+ bl_0_40 br_0_40 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c40
*+ bl_0_40 br_0_40 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c40
*+ bl_0_40 br_0_40 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c40
*+ bl_0_40 br_0_40 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c40
*+ bl_0_40 br_0_40 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c40
*+ bl_0_40 br_0_40 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c40
*+ bl_0_40 br_0_40 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c40
*+ bl_0_40 br_0_40 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c40
*+ bl_0_40 br_0_40 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c40
*+ bl_0_40 br_0_40 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c40
*+ bl_0_40 br_0_40 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c40
*+ bl_0_40 br_0_40 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c40
*+ bl_0_40 br_0_40 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c40
*+ bl_0_40 br_0_40 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c40
*+ bl_0_40 br_0_40 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c40
*+ bl_0_40 br_0_40 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c40
*+ bl_0_40 br_0_40 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c40
*+ bl_0_40 br_0_40 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c40
*+ bl_0_40 br_0_40 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c40
*+ bl_0_40 br_0_40 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c40
*+ bl_0_40 br_0_40 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c40
*+ bl_0_40 br_0_40 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c40
*+ bl_0_40 br_0_40 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c40
*+ bl_0_40 br_0_40 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c40
*+ bl_0_40 br_0_40 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c40
*+ bl_0_40 br_0_40 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c40
*+ bl_0_40 br_0_40 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c40
*+ bl_0_40 br_0_40 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c40
*+ bl_0_40 br_0_40 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c40
*+ bl_0_40 br_0_40 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c40
*+ bl_0_40 br_0_40 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c40
*+ bl_0_40 br_0_40 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c40
*+ bl_0_40 br_0_40 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c40
*+ bl_0_40 br_0_40 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c40
*+ bl_0_40 br_0_40 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c40
*+ bl_0_40 br_0_40 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c40
*+ bl_0_40 br_0_40 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c40
*+ bl_0_40 br_0_40 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c40
*+ bl_0_40 br_0_40 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c40
*+ bl_0_40 br_0_40 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c40
*+ bl_0_40 br_0_40 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c40
*+ bl_0_40 br_0_40 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c40
*+ bl_0_40 br_0_40 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c40
*+ bl_0_40 br_0_40 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c40
*+ bl_0_40 br_0_40 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c40
*+ bl_0_40 br_0_40 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c40
*+ bl_0_40 br_0_40 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c40
*+ bl_0_40 br_0_40 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c40
*+ bl_0_40 br_0_40 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c40
*+ bl_0_40 br_0_40 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c40
*+ bl_0_40 br_0_40 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c40
+ bl_0_40 br_0_40 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c41
+ bl_0_41 br_0_41 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c41
*+ bl_0_41 br_0_41 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c41
*+ bl_0_41 br_0_41 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c41
*+ bl_0_41 br_0_41 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c41
*+ bl_0_41 br_0_41 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c41
*+ bl_0_41 br_0_41 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c41
*+ bl_0_41 br_0_41 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c41
*+ bl_0_41 br_0_41 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c41
*+ bl_0_41 br_0_41 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c41
*+ bl_0_41 br_0_41 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c41
*+ bl_0_41 br_0_41 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c41
*+ bl_0_41 br_0_41 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c41
*+ bl_0_41 br_0_41 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c41
*+ bl_0_41 br_0_41 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c41
*+ bl_0_41 br_0_41 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c41
*+ bl_0_41 br_0_41 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c41
*+ bl_0_41 br_0_41 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c41
*+ bl_0_41 br_0_41 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c41
*+ bl_0_41 br_0_41 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c41
*+ bl_0_41 br_0_41 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c41
*+ bl_0_41 br_0_41 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c41
*+ bl_0_41 br_0_41 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c41
*+ bl_0_41 br_0_41 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c41
*+ bl_0_41 br_0_41 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c41
*+ bl_0_41 br_0_41 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c41
*+ bl_0_41 br_0_41 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c41
*+ bl_0_41 br_0_41 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c41
*+ bl_0_41 br_0_41 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c41
*+ bl_0_41 br_0_41 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c41
*+ bl_0_41 br_0_41 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c41
*+ bl_0_41 br_0_41 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c41
*+ bl_0_41 br_0_41 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c41
*+ bl_0_41 br_0_41 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c41
*+ bl_0_41 br_0_41 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c41
*+ bl_0_41 br_0_41 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c41
*+ bl_0_41 br_0_41 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c41
*+ bl_0_41 br_0_41 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c41
*+ bl_0_41 br_0_41 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c41
*+ bl_0_41 br_0_41 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c41
*+ bl_0_41 br_0_41 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c41
*+ bl_0_41 br_0_41 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c41
*+ bl_0_41 br_0_41 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c41
*+ bl_0_41 br_0_41 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c41
*+ bl_0_41 br_0_41 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c41
*+ bl_0_41 br_0_41 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c41
*+ bl_0_41 br_0_41 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c41
*+ bl_0_41 br_0_41 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c41
*+ bl_0_41 br_0_41 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c41
*+ bl_0_41 br_0_41 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c41
*+ bl_0_41 br_0_41 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c41
*+ bl_0_41 br_0_41 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c41
*+ bl_0_41 br_0_41 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c41
*+ bl_0_41 br_0_41 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c41
*+ bl_0_41 br_0_41 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c41
*+ bl_0_41 br_0_41 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c41
*+ bl_0_41 br_0_41 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c41
*+ bl_0_41 br_0_41 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c41
*+ bl_0_41 br_0_41 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c41
*+ bl_0_41 br_0_41 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c41
*+ bl_0_41 br_0_41 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c41
*+ bl_0_41 br_0_41 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c41
*+ bl_0_41 br_0_41 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c41
*+ bl_0_41 br_0_41 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c41
*+ bl_0_41 br_0_41 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c41
*+ bl_0_41 br_0_41 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c41
*+ bl_0_41 br_0_41 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c41
*+ bl_0_41 br_0_41 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c41
*+ bl_0_41 br_0_41 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c41
*+ bl_0_41 br_0_41 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c41
*+ bl_0_41 br_0_41 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c41
*+ bl_0_41 br_0_41 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c41
*+ bl_0_41 br_0_41 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c41
*+ bl_0_41 br_0_41 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c41
*+ bl_0_41 br_0_41 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c41
*+ bl_0_41 br_0_41 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c41
*+ bl_0_41 br_0_41 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c41
*+ bl_0_41 br_0_41 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c41
*+ bl_0_41 br_0_41 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c41
*+ bl_0_41 br_0_41 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c41
*+ bl_0_41 br_0_41 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c41
*+ bl_0_41 br_0_41 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c41
*+ bl_0_41 br_0_41 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c41
*+ bl_0_41 br_0_41 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c41
*+ bl_0_41 br_0_41 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c41
*+ bl_0_41 br_0_41 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c41
*+ bl_0_41 br_0_41 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c41
*+ bl_0_41 br_0_41 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c41
*+ bl_0_41 br_0_41 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c41
*+ bl_0_41 br_0_41 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c41
*+ bl_0_41 br_0_41 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c41
*+ bl_0_41 br_0_41 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c41
*+ bl_0_41 br_0_41 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c41
*+ bl_0_41 br_0_41 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c41
*+ bl_0_41 br_0_41 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c41
*+ bl_0_41 br_0_41 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c41
*+ bl_0_41 br_0_41 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c41
*+ bl_0_41 br_0_41 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c41
*+ bl_0_41 br_0_41 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c41
*+ bl_0_41 br_0_41 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c41
*+ bl_0_41 br_0_41 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c41
*+ bl_0_41 br_0_41 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c41
*+ bl_0_41 br_0_41 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c41
*+ bl_0_41 br_0_41 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c41
*+ bl_0_41 br_0_41 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c41
*+ bl_0_41 br_0_41 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c41
*+ bl_0_41 br_0_41 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c41
*+ bl_0_41 br_0_41 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c41
*+ bl_0_41 br_0_41 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c41
*+ bl_0_41 br_0_41 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c41
*+ bl_0_41 br_0_41 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c41
*+ bl_0_41 br_0_41 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c41
*+ bl_0_41 br_0_41 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c41
*+ bl_0_41 br_0_41 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c41
*+ bl_0_41 br_0_41 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c41
*+ bl_0_41 br_0_41 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c41
*+ bl_0_41 br_0_41 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c41
*+ bl_0_41 br_0_41 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c41
*+ bl_0_41 br_0_41 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c41
*+ bl_0_41 br_0_41 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c41
*+ bl_0_41 br_0_41 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c41
*+ bl_0_41 br_0_41 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c41
*+ bl_0_41 br_0_41 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c41
*+ bl_0_41 br_0_41 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c41
*+ bl_0_41 br_0_41 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c41
*+ bl_0_41 br_0_41 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c41
*+ bl_0_41 br_0_41 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c41
*+ bl_0_41 br_0_41 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c41
+ bl_0_41 br_0_41 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c42
+ bl_0_42 br_0_42 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c42
*+ bl_0_42 br_0_42 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c42
*+ bl_0_42 br_0_42 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c42
*+ bl_0_42 br_0_42 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c42
*+ bl_0_42 br_0_42 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c42
*+ bl_0_42 br_0_42 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c42
*+ bl_0_42 br_0_42 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c42
*+ bl_0_42 br_0_42 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c42
*+ bl_0_42 br_0_42 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c42
*+ bl_0_42 br_0_42 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c42
*+ bl_0_42 br_0_42 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c42
*+ bl_0_42 br_0_42 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c42
*+ bl_0_42 br_0_42 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c42
*+ bl_0_42 br_0_42 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c42
*+ bl_0_42 br_0_42 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c42
*+ bl_0_42 br_0_42 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c42
*+ bl_0_42 br_0_42 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c42
*+ bl_0_42 br_0_42 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c42
*+ bl_0_42 br_0_42 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c42
*+ bl_0_42 br_0_42 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c42
*+ bl_0_42 br_0_42 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c42
*+ bl_0_42 br_0_42 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c42
*+ bl_0_42 br_0_42 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c42
*+ bl_0_42 br_0_42 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c42
*+ bl_0_42 br_0_42 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c42
*+ bl_0_42 br_0_42 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c42
*+ bl_0_42 br_0_42 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c42
*+ bl_0_42 br_0_42 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c42
*+ bl_0_42 br_0_42 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c42
*+ bl_0_42 br_0_42 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c42
*+ bl_0_42 br_0_42 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c42
*+ bl_0_42 br_0_42 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c42
*+ bl_0_42 br_0_42 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c42
*+ bl_0_42 br_0_42 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c42
*+ bl_0_42 br_0_42 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c42
*+ bl_0_42 br_0_42 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c42
*+ bl_0_42 br_0_42 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c42
*+ bl_0_42 br_0_42 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c42
*+ bl_0_42 br_0_42 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c42
*+ bl_0_42 br_0_42 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c42
*+ bl_0_42 br_0_42 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c42
*+ bl_0_42 br_0_42 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c42
*+ bl_0_42 br_0_42 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c42
*+ bl_0_42 br_0_42 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c42
*+ bl_0_42 br_0_42 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c42
*+ bl_0_42 br_0_42 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c42
*+ bl_0_42 br_0_42 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c42
*+ bl_0_42 br_0_42 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c42
*+ bl_0_42 br_0_42 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c42
*+ bl_0_42 br_0_42 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c42
*+ bl_0_42 br_0_42 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c42
*+ bl_0_42 br_0_42 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c42
*+ bl_0_42 br_0_42 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c42
*+ bl_0_42 br_0_42 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c42
*+ bl_0_42 br_0_42 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c42
*+ bl_0_42 br_0_42 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c42
*+ bl_0_42 br_0_42 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c42
*+ bl_0_42 br_0_42 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c42
*+ bl_0_42 br_0_42 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c42
*+ bl_0_42 br_0_42 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c42
*+ bl_0_42 br_0_42 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c42
*+ bl_0_42 br_0_42 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c42
*+ bl_0_42 br_0_42 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c42
*+ bl_0_42 br_0_42 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c42
*+ bl_0_42 br_0_42 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c42
*+ bl_0_42 br_0_42 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c42
*+ bl_0_42 br_0_42 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c42
*+ bl_0_42 br_0_42 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c42
*+ bl_0_42 br_0_42 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c42
*+ bl_0_42 br_0_42 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c42
*+ bl_0_42 br_0_42 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c42
*+ bl_0_42 br_0_42 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c42
*+ bl_0_42 br_0_42 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c42
*+ bl_0_42 br_0_42 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c42
*+ bl_0_42 br_0_42 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c42
*+ bl_0_42 br_0_42 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c42
*+ bl_0_42 br_0_42 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c42
*+ bl_0_42 br_0_42 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c42
*+ bl_0_42 br_0_42 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c42
*+ bl_0_42 br_0_42 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c42
*+ bl_0_42 br_0_42 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c42
*+ bl_0_42 br_0_42 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c42
*+ bl_0_42 br_0_42 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c42
*+ bl_0_42 br_0_42 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c42
*+ bl_0_42 br_0_42 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c42
*+ bl_0_42 br_0_42 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c42
*+ bl_0_42 br_0_42 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c42
*+ bl_0_42 br_0_42 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c42
*+ bl_0_42 br_0_42 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c42
*+ bl_0_42 br_0_42 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c42
*+ bl_0_42 br_0_42 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c42
*+ bl_0_42 br_0_42 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c42
*+ bl_0_42 br_0_42 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c42
*+ bl_0_42 br_0_42 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c42
*+ bl_0_42 br_0_42 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c42
*+ bl_0_42 br_0_42 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c42
*+ bl_0_42 br_0_42 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c42
*+ bl_0_42 br_0_42 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c42
*+ bl_0_42 br_0_42 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c42
*+ bl_0_42 br_0_42 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c42
*+ bl_0_42 br_0_42 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c42
*+ bl_0_42 br_0_42 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c42
*+ bl_0_42 br_0_42 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c42
*+ bl_0_42 br_0_42 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c42
*+ bl_0_42 br_0_42 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c42
*+ bl_0_42 br_0_42 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c42
*+ bl_0_42 br_0_42 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c42
*+ bl_0_42 br_0_42 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c42
*+ bl_0_42 br_0_42 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c42
*+ bl_0_42 br_0_42 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c42
*+ bl_0_42 br_0_42 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c42
*+ bl_0_42 br_0_42 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c42
*+ bl_0_42 br_0_42 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c42
*+ bl_0_42 br_0_42 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c42
*+ bl_0_42 br_0_42 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c42
*+ bl_0_42 br_0_42 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c42
*+ bl_0_42 br_0_42 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c42
*+ bl_0_42 br_0_42 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c42
*+ bl_0_42 br_0_42 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c42
*+ bl_0_42 br_0_42 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c42
*+ bl_0_42 br_0_42 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c42
*+ bl_0_42 br_0_42 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c42
*+ bl_0_42 br_0_42 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c42
*+ bl_0_42 br_0_42 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c42
*+ bl_0_42 br_0_42 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c42
*+ bl_0_42 br_0_42 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c42
*+ bl_0_42 br_0_42 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c42
+ bl_0_42 br_0_42 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c43
+ bl_0_43 br_0_43 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c43
*+ bl_0_43 br_0_43 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c43
*+ bl_0_43 br_0_43 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c43
*+ bl_0_43 br_0_43 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c43
*+ bl_0_43 br_0_43 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c43
*+ bl_0_43 br_0_43 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c43
*+ bl_0_43 br_0_43 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c43
*+ bl_0_43 br_0_43 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c43
*+ bl_0_43 br_0_43 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c43
*+ bl_0_43 br_0_43 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c43
*+ bl_0_43 br_0_43 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c43
*+ bl_0_43 br_0_43 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c43
*+ bl_0_43 br_0_43 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c43
*+ bl_0_43 br_0_43 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c43
*+ bl_0_43 br_0_43 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c43
*+ bl_0_43 br_0_43 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c43
*+ bl_0_43 br_0_43 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c43
*+ bl_0_43 br_0_43 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c43
*+ bl_0_43 br_0_43 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c43
*+ bl_0_43 br_0_43 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c43
*+ bl_0_43 br_0_43 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c43
*+ bl_0_43 br_0_43 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c43
*+ bl_0_43 br_0_43 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c43
*+ bl_0_43 br_0_43 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c43
*+ bl_0_43 br_0_43 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c43
*+ bl_0_43 br_0_43 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c43
*+ bl_0_43 br_0_43 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c43
*+ bl_0_43 br_0_43 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c43
*+ bl_0_43 br_0_43 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c43
*+ bl_0_43 br_0_43 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c43
*+ bl_0_43 br_0_43 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c43
*+ bl_0_43 br_0_43 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c43
*+ bl_0_43 br_0_43 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c43
*+ bl_0_43 br_0_43 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c43
*+ bl_0_43 br_0_43 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c43
*+ bl_0_43 br_0_43 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c43
*+ bl_0_43 br_0_43 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c43
*+ bl_0_43 br_0_43 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c43
*+ bl_0_43 br_0_43 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c43
*+ bl_0_43 br_0_43 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c43
*+ bl_0_43 br_0_43 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c43
*+ bl_0_43 br_0_43 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c43
*+ bl_0_43 br_0_43 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c43
*+ bl_0_43 br_0_43 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c43
*+ bl_0_43 br_0_43 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c43
*+ bl_0_43 br_0_43 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c43
*+ bl_0_43 br_0_43 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c43
*+ bl_0_43 br_0_43 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c43
*+ bl_0_43 br_0_43 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c43
*+ bl_0_43 br_0_43 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c43
*+ bl_0_43 br_0_43 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c43
*+ bl_0_43 br_0_43 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c43
*+ bl_0_43 br_0_43 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c43
*+ bl_0_43 br_0_43 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c43
*+ bl_0_43 br_0_43 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c43
*+ bl_0_43 br_0_43 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c43
*+ bl_0_43 br_0_43 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c43
*+ bl_0_43 br_0_43 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c43
*+ bl_0_43 br_0_43 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c43
*+ bl_0_43 br_0_43 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c43
*+ bl_0_43 br_0_43 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c43
*+ bl_0_43 br_0_43 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c43
*+ bl_0_43 br_0_43 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c43
*+ bl_0_43 br_0_43 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c43
*+ bl_0_43 br_0_43 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c43
*+ bl_0_43 br_0_43 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c43
*+ bl_0_43 br_0_43 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c43
*+ bl_0_43 br_0_43 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c43
*+ bl_0_43 br_0_43 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c43
*+ bl_0_43 br_0_43 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c43
*+ bl_0_43 br_0_43 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c43
*+ bl_0_43 br_0_43 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c43
*+ bl_0_43 br_0_43 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c43
*+ bl_0_43 br_0_43 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c43
*+ bl_0_43 br_0_43 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c43
*+ bl_0_43 br_0_43 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c43
*+ bl_0_43 br_0_43 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c43
*+ bl_0_43 br_0_43 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c43
*+ bl_0_43 br_0_43 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c43
*+ bl_0_43 br_0_43 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c43
*+ bl_0_43 br_0_43 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c43
*+ bl_0_43 br_0_43 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c43
*+ bl_0_43 br_0_43 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c43
*+ bl_0_43 br_0_43 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c43
*+ bl_0_43 br_0_43 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c43
*+ bl_0_43 br_0_43 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c43
*+ bl_0_43 br_0_43 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c43
*+ bl_0_43 br_0_43 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c43
*+ bl_0_43 br_0_43 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c43
*+ bl_0_43 br_0_43 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c43
*+ bl_0_43 br_0_43 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c43
*+ bl_0_43 br_0_43 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c43
*+ bl_0_43 br_0_43 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c43
*+ bl_0_43 br_0_43 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c43
*+ bl_0_43 br_0_43 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c43
*+ bl_0_43 br_0_43 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c43
*+ bl_0_43 br_0_43 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c43
*+ bl_0_43 br_0_43 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c43
*+ bl_0_43 br_0_43 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c43
*+ bl_0_43 br_0_43 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c43
*+ bl_0_43 br_0_43 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c43
*+ bl_0_43 br_0_43 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c43
*+ bl_0_43 br_0_43 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c43
*+ bl_0_43 br_0_43 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c43
*+ bl_0_43 br_0_43 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c43
*+ bl_0_43 br_0_43 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c43
*+ bl_0_43 br_0_43 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c43
*+ bl_0_43 br_0_43 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c43
*+ bl_0_43 br_0_43 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c43
*+ bl_0_43 br_0_43 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c43
*+ bl_0_43 br_0_43 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c43
*+ bl_0_43 br_0_43 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c43
*+ bl_0_43 br_0_43 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c43
*+ bl_0_43 br_0_43 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c43
*+ bl_0_43 br_0_43 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c43
*+ bl_0_43 br_0_43 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c43
*+ bl_0_43 br_0_43 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c43
*+ bl_0_43 br_0_43 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c43
*+ bl_0_43 br_0_43 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c43
*+ bl_0_43 br_0_43 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c43
*+ bl_0_43 br_0_43 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c43
*+ bl_0_43 br_0_43 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c43
*+ bl_0_43 br_0_43 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c43
*+ bl_0_43 br_0_43 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c43
*+ bl_0_43 br_0_43 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c43
*+ bl_0_43 br_0_43 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c43
*+ bl_0_43 br_0_43 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c43
+ bl_0_43 br_0_43 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c44
+ bl_0_44 br_0_44 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c44
*+ bl_0_44 br_0_44 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c44
*+ bl_0_44 br_0_44 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c44
*+ bl_0_44 br_0_44 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c44
*+ bl_0_44 br_0_44 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c44
*+ bl_0_44 br_0_44 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c44
*+ bl_0_44 br_0_44 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c44
*+ bl_0_44 br_0_44 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c44
*+ bl_0_44 br_0_44 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c44
*+ bl_0_44 br_0_44 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c44
*+ bl_0_44 br_0_44 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c44
*+ bl_0_44 br_0_44 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c44
*+ bl_0_44 br_0_44 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c44
*+ bl_0_44 br_0_44 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c44
*+ bl_0_44 br_0_44 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c44
*+ bl_0_44 br_0_44 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c44
*+ bl_0_44 br_0_44 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c44
*+ bl_0_44 br_0_44 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c44
*+ bl_0_44 br_0_44 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c44
*+ bl_0_44 br_0_44 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c44
*+ bl_0_44 br_0_44 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c44
*+ bl_0_44 br_0_44 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c44
*+ bl_0_44 br_0_44 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c44
*+ bl_0_44 br_0_44 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c44
*+ bl_0_44 br_0_44 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c44
*+ bl_0_44 br_0_44 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c44
*+ bl_0_44 br_0_44 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c44
*+ bl_0_44 br_0_44 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c44
*+ bl_0_44 br_0_44 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c44
*+ bl_0_44 br_0_44 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c44
*+ bl_0_44 br_0_44 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c44
*+ bl_0_44 br_0_44 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c44
*+ bl_0_44 br_0_44 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c44
*+ bl_0_44 br_0_44 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c44
*+ bl_0_44 br_0_44 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c44
*+ bl_0_44 br_0_44 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c44
*+ bl_0_44 br_0_44 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c44
*+ bl_0_44 br_0_44 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c44
*+ bl_0_44 br_0_44 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c44
*+ bl_0_44 br_0_44 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c44
*+ bl_0_44 br_0_44 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c44
*+ bl_0_44 br_0_44 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c44
*+ bl_0_44 br_0_44 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c44
*+ bl_0_44 br_0_44 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c44
*+ bl_0_44 br_0_44 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c44
*+ bl_0_44 br_0_44 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c44
*+ bl_0_44 br_0_44 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c44
*+ bl_0_44 br_0_44 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c44
*+ bl_0_44 br_0_44 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c44
*+ bl_0_44 br_0_44 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c44
*+ bl_0_44 br_0_44 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c44
*+ bl_0_44 br_0_44 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c44
*+ bl_0_44 br_0_44 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c44
*+ bl_0_44 br_0_44 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c44
*+ bl_0_44 br_0_44 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c44
*+ bl_0_44 br_0_44 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c44
*+ bl_0_44 br_0_44 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c44
*+ bl_0_44 br_0_44 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c44
*+ bl_0_44 br_0_44 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c44
*+ bl_0_44 br_0_44 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c44
*+ bl_0_44 br_0_44 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c44
*+ bl_0_44 br_0_44 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c44
*+ bl_0_44 br_0_44 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c44
*+ bl_0_44 br_0_44 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c44
*+ bl_0_44 br_0_44 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c44
*+ bl_0_44 br_0_44 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c44
*+ bl_0_44 br_0_44 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c44
*+ bl_0_44 br_0_44 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c44
*+ bl_0_44 br_0_44 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c44
*+ bl_0_44 br_0_44 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c44
*+ bl_0_44 br_0_44 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c44
*+ bl_0_44 br_0_44 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c44
*+ bl_0_44 br_0_44 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c44
*+ bl_0_44 br_0_44 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c44
*+ bl_0_44 br_0_44 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c44
*+ bl_0_44 br_0_44 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c44
*+ bl_0_44 br_0_44 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c44
*+ bl_0_44 br_0_44 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c44
*+ bl_0_44 br_0_44 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c44
*+ bl_0_44 br_0_44 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c44
*+ bl_0_44 br_0_44 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c44
*+ bl_0_44 br_0_44 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c44
*+ bl_0_44 br_0_44 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c44
*+ bl_0_44 br_0_44 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c44
*+ bl_0_44 br_0_44 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c44
*+ bl_0_44 br_0_44 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c44
*+ bl_0_44 br_0_44 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c44
*+ bl_0_44 br_0_44 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c44
*+ bl_0_44 br_0_44 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c44
*+ bl_0_44 br_0_44 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c44
*+ bl_0_44 br_0_44 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c44
*+ bl_0_44 br_0_44 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c44
*+ bl_0_44 br_0_44 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c44
*+ bl_0_44 br_0_44 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c44
*+ bl_0_44 br_0_44 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c44
*+ bl_0_44 br_0_44 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c44
*+ bl_0_44 br_0_44 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c44
*+ bl_0_44 br_0_44 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c44
*+ bl_0_44 br_0_44 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c44
*+ bl_0_44 br_0_44 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c44
*+ bl_0_44 br_0_44 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c44
*+ bl_0_44 br_0_44 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c44
*+ bl_0_44 br_0_44 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c44
*+ bl_0_44 br_0_44 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c44
*+ bl_0_44 br_0_44 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c44
*+ bl_0_44 br_0_44 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c44
*+ bl_0_44 br_0_44 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c44
*+ bl_0_44 br_0_44 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c44
*+ bl_0_44 br_0_44 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c44
*+ bl_0_44 br_0_44 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c44
*+ bl_0_44 br_0_44 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c44
*+ bl_0_44 br_0_44 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c44
*+ bl_0_44 br_0_44 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c44
*+ bl_0_44 br_0_44 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c44
*+ bl_0_44 br_0_44 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c44
*+ bl_0_44 br_0_44 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c44
*+ bl_0_44 br_0_44 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c44
*+ bl_0_44 br_0_44 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c44
*+ bl_0_44 br_0_44 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c44
*+ bl_0_44 br_0_44 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c44
*+ bl_0_44 br_0_44 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c44
*+ bl_0_44 br_0_44 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c44
*+ bl_0_44 br_0_44 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c44
*+ bl_0_44 br_0_44 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c44
*+ bl_0_44 br_0_44 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c44
*+ bl_0_44 br_0_44 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c44
*+ bl_0_44 br_0_44 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c44
+ bl_0_44 br_0_44 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c45
+ bl_0_45 br_0_45 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c45
*+ bl_0_45 br_0_45 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c45
*+ bl_0_45 br_0_45 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c45
*+ bl_0_45 br_0_45 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c45
*+ bl_0_45 br_0_45 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c45
*+ bl_0_45 br_0_45 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c45
*+ bl_0_45 br_0_45 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c45
*+ bl_0_45 br_0_45 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c45
*+ bl_0_45 br_0_45 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c45
*+ bl_0_45 br_0_45 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c45
*+ bl_0_45 br_0_45 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c45
*+ bl_0_45 br_0_45 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c45
*+ bl_0_45 br_0_45 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c45
*+ bl_0_45 br_0_45 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c45
*+ bl_0_45 br_0_45 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c45
*+ bl_0_45 br_0_45 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c45
*+ bl_0_45 br_0_45 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c45
*+ bl_0_45 br_0_45 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c45
*+ bl_0_45 br_0_45 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c45
*+ bl_0_45 br_0_45 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c45
*+ bl_0_45 br_0_45 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c45
*+ bl_0_45 br_0_45 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c45
*+ bl_0_45 br_0_45 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c45
*+ bl_0_45 br_0_45 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c45
*+ bl_0_45 br_0_45 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c45
*+ bl_0_45 br_0_45 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c45
*+ bl_0_45 br_0_45 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c45
*+ bl_0_45 br_0_45 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c45
*+ bl_0_45 br_0_45 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c45
*+ bl_0_45 br_0_45 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c45
*+ bl_0_45 br_0_45 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c45
*+ bl_0_45 br_0_45 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c45
*+ bl_0_45 br_0_45 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c45
*+ bl_0_45 br_0_45 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c45
*+ bl_0_45 br_0_45 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c45
*+ bl_0_45 br_0_45 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c45
*+ bl_0_45 br_0_45 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c45
*+ bl_0_45 br_0_45 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c45
*+ bl_0_45 br_0_45 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c45
*+ bl_0_45 br_0_45 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c45
*+ bl_0_45 br_0_45 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c45
*+ bl_0_45 br_0_45 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c45
*+ bl_0_45 br_0_45 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c45
*+ bl_0_45 br_0_45 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c45
*+ bl_0_45 br_0_45 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c45
*+ bl_0_45 br_0_45 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c45
*+ bl_0_45 br_0_45 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c45
*+ bl_0_45 br_0_45 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c45
*+ bl_0_45 br_0_45 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c45
*+ bl_0_45 br_0_45 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c45
*+ bl_0_45 br_0_45 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c45
*+ bl_0_45 br_0_45 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c45
*+ bl_0_45 br_0_45 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c45
*+ bl_0_45 br_0_45 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c45
*+ bl_0_45 br_0_45 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c45
*+ bl_0_45 br_0_45 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c45
*+ bl_0_45 br_0_45 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c45
*+ bl_0_45 br_0_45 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c45
*+ bl_0_45 br_0_45 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c45
*+ bl_0_45 br_0_45 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c45
*+ bl_0_45 br_0_45 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c45
*+ bl_0_45 br_0_45 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c45
*+ bl_0_45 br_0_45 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c45
*+ bl_0_45 br_0_45 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c45
*+ bl_0_45 br_0_45 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c45
*+ bl_0_45 br_0_45 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c45
*+ bl_0_45 br_0_45 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c45
*+ bl_0_45 br_0_45 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c45
*+ bl_0_45 br_0_45 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c45
*+ bl_0_45 br_0_45 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c45
*+ bl_0_45 br_0_45 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c45
*+ bl_0_45 br_0_45 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c45
*+ bl_0_45 br_0_45 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c45
*+ bl_0_45 br_0_45 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c45
*+ bl_0_45 br_0_45 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c45
*+ bl_0_45 br_0_45 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c45
*+ bl_0_45 br_0_45 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c45
*+ bl_0_45 br_0_45 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c45
*+ bl_0_45 br_0_45 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c45
*+ bl_0_45 br_0_45 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c45
*+ bl_0_45 br_0_45 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c45
*+ bl_0_45 br_0_45 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c45
*+ bl_0_45 br_0_45 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c45
*+ bl_0_45 br_0_45 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c45
*+ bl_0_45 br_0_45 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c45
*+ bl_0_45 br_0_45 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c45
*+ bl_0_45 br_0_45 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c45
*+ bl_0_45 br_0_45 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c45
*+ bl_0_45 br_0_45 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c45
*+ bl_0_45 br_0_45 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c45
*+ bl_0_45 br_0_45 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c45
*+ bl_0_45 br_0_45 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c45
*+ bl_0_45 br_0_45 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c45
*+ bl_0_45 br_0_45 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c45
*+ bl_0_45 br_0_45 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c45
*+ bl_0_45 br_0_45 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c45
*+ bl_0_45 br_0_45 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c45
*+ bl_0_45 br_0_45 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c45
*+ bl_0_45 br_0_45 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c45
*+ bl_0_45 br_0_45 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c45
*+ bl_0_45 br_0_45 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c45
*+ bl_0_45 br_0_45 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c45
*+ bl_0_45 br_0_45 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c45
*+ bl_0_45 br_0_45 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c45
*+ bl_0_45 br_0_45 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c45
*+ bl_0_45 br_0_45 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c45
*+ bl_0_45 br_0_45 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c45
*+ bl_0_45 br_0_45 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c45
*+ bl_0_45 br_0_45 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c45
*+ bl_0_45 br_0_45 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c45
*+ bl_0_45 br_0_45 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c45
*+ bl_0_45 br_0_45 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c45
*+ bl_0_45 br_0_45 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c45
*+ bl_0_45 br_0_45 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c45
*+ bl_0_45 br_0_45 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c45
*+ bl_0_45 br_0_45 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c45
*+ bl_0_45 br_0_45 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c45
*+ bl_0_45 br_0_45 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c45
*+ bl_0_45 br_0_45 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c45
*+ bl_0_45 br_0_45 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c45
*+ bl_0_45 br_0_45 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c45
*+ bl_0_45 br_0_45 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c45
*+ bl_0_45 br_0_45 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c45
*+ bl_0_45 br_0_45 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c45
*+ bl_0_45 br_0_45 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c45
*+ bl_0_45 br_0_45 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c45
*+ bl_0_45 br_0_45 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c45
+ bl_0_45 br_0_45 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c46
+ bl_0_46 br_0_46 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c46
*+ bl_0_46 br_0_46 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c46
*+ bl_0_46 br_0_46 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c46
*+ bl_0_46 br_0_46 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c46
*+ bl_0_46 br_0_46 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c46
*+ bl_0_46 br_0_46 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c46
*+ bl_0_46 br_0_46 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c46
*+ bl_0_46 br_0_46 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c46
*+ bl_0_46 br_0_46 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c46
*+ bl_0_46 br_0_46 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c46
*+ bl_0_46 br_0_46 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c46
*+ bl_0_46 br_0_46 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c46
*+ bl_0_46 br_0_46 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c46
*+ bl_0_46 br_0_46 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c46
*+ bl_0_46 br_0_46 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c46
*+ bl_0_46 br_0_46 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c46
*+ bl_0_46 br_0_46 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c46
*+ bl_0_46 br_0_46 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c46
*+ bl_0_46 br_0_46 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c46
*+ bl_0_46 br_0_46 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c46
*+ bl_0_46 br_0_46 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c46
*+ bl_0_46 br_0_46 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c46
*+ bl_0_46 br_0_46 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c46
*+ bl_0_46 br_0_46 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c46
*+ bl_0_46 br_0_46 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c46
*+ bl_0_46 br_0_46 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c46
*+ bl_0_46 br_0_46 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c46
*+ bl_0_46 br_0_46 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c46
*+ bl_0_46 br_0_46 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c46
*+ bl_0_46 br_0_46 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c46
*+ bl_0_46 br_0_46 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c46
*+ bl_0_46 br_0_46 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c46
*+ bl_0_46 br_0_46 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c46
*+ bl_0_46 br_0_46 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c46
*+ bl_0_46 br_0_46 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c46
*+ bl_0_46 br_0_46 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c46
*+ bl_0_46 br_0_46 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c46
*+ bl_0_46 br_0_46 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c46
*+ bl_0_46 br_0_46 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c46
*+ bl_0_46 br_0_46 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c46
*+ bl_0_46 br_0_46 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c46
*+ bl_0_46 br_0_46 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c46
*+ bl_0_46 br_0_46 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c46
*+ bl_0_46 br_0_46 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c46
*+ bl_0_46 br_0_46 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c46
*+ bl_0_46 br_0_46 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c46
*+ bl_0_46 br_0_46 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c46
*+ bl_0_46 br_0_46 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c46
*+ bl_0_46 br_0_46 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c46
*+ bl_0_46 br_0_46 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c46
*+ bl_0_46 br_0_46 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c46
*+ bl_0_46 br_0_46 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c46
*+ bl_0_46 br_0_46 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c46
*+ bl_0_46 br_0_46 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c46
*+ bl_0_46 br_0_46 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c46
*+ bl_0_46 br_0_46 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c46
*+ bl_0_46 br_0_46 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c46
*+ bl_0_46 br_0_46 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c46
*+ bl_0_46 br_0_46 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c46
*+ bl_0_46 br_0_46 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c46
*+ bl_0_46 br_0_46 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c46
*+ bl_0_46 br_0_46 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c46
*+ bl_0_46 br_0_46 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c46
*+ bl_0_46 br_0_46 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c46
*+ bl_0_46 br_0_46 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c46
*+ bl_0_46 br_0_46 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c46
*+ bl_0_46 br_0_46 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c46
*+ bl_0_46 br_0_46 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c46
*+ bl_0_46 br_0_46 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c46
*+ bl_0_46 br_0_46 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c46
*+ bl_0_46 br_0_46 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c46
*+ bl_0_46 br_0_46 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c46
*+ bl_0_46 br_0_46 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c46
*+ bl_0_46 br_0_46 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c46
*+ bl_0_46 br_0_46 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c46
*+ bl_0_46 br_0_46 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c46
*+ bl_0_46 br_0_46 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c46
*+ bl_0_46 br_0_46 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c46
*+ bl_0_46 br_0_46 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c46
*+ bl_0_46 br_0_46 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c46
*+ bl_0_46 br_0_46 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c46
*+ bl_0_46 br_0_46 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c46
*+ bl_0_46 br_0_46 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c46
*+ bl_0_46 br_0_46 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c46
*+ bl_0_46 br_0_46 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c46
*+ bl_0_46 br_0_46 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c46
*+ bl_0_46 br_0_46 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c46
*+ bl_0_46 br_0_46 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c46
*+ bl_0_46 br_0_46 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c46
*+ bl_0_46 br_0_46 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c46
*+ bl_0_46 br_0_46 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c46
*+ bl_0_46 br_0_46 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c46
*+ bl_0_46 br_0_46 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c46
*+ bl_0_46 br_0_46 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c46
*+ bl_0_46 br_0_46 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c46
*+ bl_0_46 br_0_46 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c46
*+ bl_0_46 br_0_46 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c46
*+ bl_0_46 br_0_46 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c46
*+ bl_0_46 br_0_46 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c46
*+ bl_0_46 br_0_46 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c46
*+ bl_0_46 br_0_46 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c46
*+ bl_0_46 br_0_46 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c46
*+ bl_0_46 br_0_46 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c46
*+ bl_0_46 br_0_46 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c46
*+ bl_0_46 br_0_46 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c46
*+ bl_0_46 br_0_46 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c46
*+ bl_0_46 br_0_46 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c46
*+ bl_0_46 br_0_46 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c46
*+ bl_0_46 br_0_46 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c46
*+ bl_0_46 br_0_46 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c46
*+ bl_0_46 br_0_46 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c46
*+ bl_0_46 br_0_46 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c46
*+ bl_0_46 br_0_46 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c46
*+ bl_0_46 br_0_46 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c46
*+ bl_0_46 br_0_46 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c46
*+ bl_0_46 br_0_46 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c46
*+ bl_0_46 br_0_46 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c46
*+ bl_0_46 br_0_46 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c46
*+ bl_0_46 br_0_46 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c46
*+ bl_0_46 br_0_46 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c46
*+ bl_0_46 br_0_46 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c46
*+ bl_0_46 br_0_46 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c46
*+ bl_0_46 br_0_46 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c46
*+ bl_0_46 br_0_46 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c46
*+ bl_0_46 br_0_46 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c46
*+ bl_0_46 br_0_46 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c46
*+ bl_0_46 br_0_46 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c46
+ bl_0_46 br_0_46 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c47
+ bl_0_47 br_0_47 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c47
*+ bl_0_47 br_0_47 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c47
*+ bl_0_47 br_0_47 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c47
*+ bl_0_47 br_0_47 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c47
*+ bl_0_47 br_0_47 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c47
*+ bl_0_47 br_0_47 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c47
*+ bl_0_47 br_0_47 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c47
*+ bl_0_47 br_0_47 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c47
*+ bl_0_47 br_0_47 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c47
*+ bl_0_47 br_0_47 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c47
*+ bl_0_47 br_0_47 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c47
*+ bl_0_47 br_0_47 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c47
*+ bl_0_47 br_0_47 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c47
*+ bl_0_47 br_0_47 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c47
*+ bl_0_47 br_0_47 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c47
*+ bl_0_47 br_0_47 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c47
*+ bl_0_47 br_0_47 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c47
*+ bl_0_47 br_0_47 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c47
*+ bl_0_47 br_0_47 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c47
*+ bl_0_47 br_0_47 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c47
*+ bl_0_47 br_0_47 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c47
*+ bl_0_47 br_0_47 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c47
*+ bl_0_47 br_0_47 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c47
*+ bl_0_47 br_0_47 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c47
*+ bl_0_47 br_0_47 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c47
*+ bl_0_47 br_0_47 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c47
*+ bl_0_47 br_0_47 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c47
*+ bl_0_47 br_0_47 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c47
*+ bl_0_47 br_0_47 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c47
*+ bl_0_47 br_0_47 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c47
*+ bl_0_47 br_0_47 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c47
*+ bl_0_47 br_0_47 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c47
*+ bl_0_47 br_0_47 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c47
*+ bl_0_47 br_0_47 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c47
*+ bl_0_47 br_0_47 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c47
*+ bl_0_47 br_0_47 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c47
*+ bl_0_47 br_0_47 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c47
*+ bl_0_47 br_0_47 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c47
*+ bl_0_47 br_0_47 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c47
*+ bl_0_47 br_0_47 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c47
*+ bl_0_47 br_0_47 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c47
*+ bl_0_47 br_0_47 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c47
*+ bl_0_47 br_0_47 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c47
*+ bl_0_47 br_0_47 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c47
*+ bl_0_47 br_0_47 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c47
*+ bl_0_47 br_0_47 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c47
*+ bl_0_47 br_0_47 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c47
*+ bl_0_47 br_0_47 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c47
*+ bl_0_47 br_0_47 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c47
*+ bl_0_47 br_0_47 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c47
*+ bl_0_47 br_0_47 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c47
*+ bl_0_47 br_0_47 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c47
*+ bl_0_47 br_0_47 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c47
*+ bl_0_47 br_0_47 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c47
*+ bl_0_47 br_0_47 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c47
*+ bl_0_47 br_0_47 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c47
*+ bl_0_47 br_0_47 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c47
*+ bl_0_47 br_0_47 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c47
*+ bl_0_47 br_0_47 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c47
*+ bl_0_47 br_0_47 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c47
*+ bl_0_47 br_0_47 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c47
*+ bl_0_47 br_0_47 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c47
*+ bl_0_47 br_0_47 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c47
*+ bl_0_47 br_0_47 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c47
*+ bl_0_47 br_0_47 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c47
*+ bl_0_47 br_0_47 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c47
*+ bl_0_47 br_0_47 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c47
*+ bl_0_47 br_0_47 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c47
*+ bl_0_47 br_0_47 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c47
*+ bl_0_47 br_0_47 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c47
*+ bl_0_47 br_0_47 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c47
*+ bl_0_47 br_0_47 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c47
*+ bl_0_47 br_0_47 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c47
*+ bl_0_47 br_0_47 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c47
*+ bl_0_47 br_0_47 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c47
*+ bl_0_47 br_0_47 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c47
*+ bl_0_47 br_0_47 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c47
*+ bl_0_47 br_0_47 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c47
*+ bl_0_47 br_0_47 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c47
*+ bl_0_47 br_0_47 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c47
*+ bl_0_47 br_0_47 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c47
*+ bl_0_47 br_0_47 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c47
*+ bl_0_47 br_0_47 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c47
*+ bl_0_47 br_0_47 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c47
*+ bl_0_47 br_0_47 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c47
*+ bl_0_47 br_0_47 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c47
*+ bl_0_47 br_0_47 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c47
*+ bl_0_47 br_0_47 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c47
*+ bl_0_47 br_0_47 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c47
*+ bl_0_47 br_0_47 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c47
*+ bl_0_47 br_0_47 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c47
*+ bl_0_47 br_0_47 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c47
*+ bl_0_47 br_0_47 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c47
*+ bl_0_47 br_0_47 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c47
*+ bl_0_47 br_0_47 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c47
*+ bl_0_47 br_0_47 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c47
*+ bl_0_47 br_0_47 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c47
*+ bl_0_47 br_0_47 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c47
*+ bl_0_47 br_0_47 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c47
*+ bl_0_47 br_0_47 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c47
*+ bl_0_47 br_0_47 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c47
*+ bl_0_47 br_0_47 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c47
*+ bl_0_47 br_0_47 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c47
*+ bl_0_47 br_0_47 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c47
*+ bl_0_47 br_0_47 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c47
*+ bl_0_47 br_0_47 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c47
*+ bl_0_47 br_0_47 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c47
*+ bl_0_47 br_0_47 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c47
*+ bl_0_47 br_0_47 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c47
*+ bl_0_47 br_0_47 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c47
*+ bl_0_47 br_0_47 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c47
*+ bl_0_47 br_0_47 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c47
*+ bl_0_47 br_0_47 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c47
*+ bl_0_47 br_0_47 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c47
*+ bl_0_47 br_0_47 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c47
*+ bl_0_47 br_0_47 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c47
*+ bl_0_47 br_0_47 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c47
*+ bl_0_47 br_0_47 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c47
*+ bl_0_47 br_0_47 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c47
*+ bl_0_47 br_0_47 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c47
*+ bl_0_47 br_0_47 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c47
*+ bl_0_47 br_0_47 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c47
*+ bl_0_47 br_0_47 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c47
*+ bl_0_47 br_0_47 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c47
*+ bl_0_47 br_0_47 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c47
*+ bl_0_47 br_0_47 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c47
*+ bl_0_47 br_0_47 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c47
+ bl_0_47 br_0_47 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c48
+ bl_0_48 br_0_48 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c48
*+ bl_0_48 br_0_48 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c48
*+ bl_0_48 br_0_48 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c48
*+ bl_0_48 br_0_48 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c48
*+ bl_0_48 br_0_48 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c48
*+ bl_0_48 br_0_48 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c48
*+ bl_0_48 br_0_48 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c48
*+ bl_0_48 br_0_48 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c48
*+ bl_0_48 br_0_48 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c48
*+ bl_0_48 br_0_48 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c48
*+ bl_0_48 br_0_48 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c48
*+ bl_0_48 br_0_48 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c48
*+ bl_0_48 br_0_48 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c48
*+ bl_0_48 br_0_48 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c48
*+ bl_0_48 br_0_48 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c48
*+ bl_0_48 br_0_48 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c48
*+ bl_0_48 br_0_48 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c48
*+ bl_0_48 br_0_48 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c48
*+ bl_0_48 br_0_48 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c48
*+ bl_0_48 br_0_48 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c48
*+ bl_0_48 br_0_48 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c48
*+ bl_0_48 br_0_48 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c48
*+ bl_0_48 br_0_48 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c48
*+ bl_0_48 br_0_48 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c48
*+ bl_0_48 br_0_48 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c48
*+ bl_0_48 br_0_48 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c48
*+ bl_0_48 br_0_48 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c48
*+ bl_0_48 br_0_48 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c48
*+ bl_0_48 br_0_48 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c48
*+ bl_0_48 br_0_48 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c48
*+ bl_0_48 br_0_48 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c48
*+ bl_0_48 br_0_48 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c48
*+ bl_0_48 br_0_48 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c48
*+ bl_0_48 br_0_48 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c48
*+ bl_0_48 br_0_48 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c48
*+ bl_0_48 br_0_48 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c48
*+ bl_0_48 br_0_48 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c48
*+ bl_0_48 br_0_48 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c48
*+ bl_0_48 br_0_48 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c48
*+ bl_0_48 br_0_48 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c48
*+ bl_0_48 br_0_48 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c48
*+ bl_0_48 br_0_48 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c48
*+ bl_0_48 br_0_48 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c48
*+ bl_0_48 br_0_48 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c48
*+ bl_0_48 br_0_48 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c48
*+ bl_0_48 br_0_48 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c48
*+ bl_0_48 br_0_48 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c48
*+ bl_0_48 br_0_48 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c48
*+ bl_0_48 br_0_48 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c48
*+ bl_0_48 br_0_48 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c48
*+ bl_0_48 br_0_48 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c48
*+ bl_0_48 br_0_48 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c48
*+ bl_0_48 br_0_48 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c48
*+ bl_0_48 br_0_48 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c48
*+ bl_0_48 br_0_48 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c48
*+ bl_0_48 br_0_48 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c48
*+ bl_0_48 br_0_48 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c48
*+ bl_0_48 br_0_48 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c48
*+ bl_0_48 br_0_48 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c48
*+ bl_0_48 br_0_48 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c48
*+ bl_0_48 br_0_48 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c48
*+ bl_0_48 br_0_48 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c48
*+ bl_0_48 br_0_48 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c48
*+ bl_0_48 br_0_48 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c48
*+ bl_0_48 br_0_48 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c48
*+ bl_0_48 br_0_48 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c48
*+ bl_0_48 br_0_48 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c48
*+ bl_0_48 br_0_48 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c48
*+ bl_0_48 br_0_48 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c48
*+ bl_0_48 br_0_48 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c48
*+ bl_0_48 br_0_48 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c48
*+ bl_0_48 br_0_48 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c48
*+ bl_0_48 br_0_48 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c48
*+ bl_0_48 br_0_48 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c48
*+ bl_0_48 br_0_48 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c48
*+ bl_0_48 br_0_48 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c48
*+ bl_0_48 br_0_48 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c48
*+ bl_0_48 br_0_48 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c48
*+ bl_0_48 br_0_48 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c48
*+ bl_0_48 br_0_48 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c48
*+ bl_0_48 br_0_48 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c48
*+ bl_0_48 br_0_48 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c48
*+ bl_0_48 br_0_48 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c48
*+ bl_0_48 br_0_48 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c48
*+ bl_0_48 br_0_48 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c48
*+ bl_0_48 br_0_48 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c48
*+ bl_0_48 br_0_48 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c48
*+ bl_0_48 br_0_48 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c48
*+ bl_0_48 br_0_48 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c48
*+ bl_0_48 br_0_48 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c48
*+ bl_0_48 br_0_48 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c48
*+ bl_0_48 br_0_48 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c48
*+ bl_0_48 br_0_48 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c48
*+ bl_0_48 br_0_48 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c48
*+ bl_0_48 br_0_48 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c48
*+ bl_0_48 br_0_48 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c48
*+ bl_0_48 br_0_48 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c48
*+ bl_0_48 br_0_48 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c48
*+ bl_0_48 br_0_48 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c48
*+ bl_0_48 br_0_48 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c48
*+ bl_0_48 br_0_48 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c48
*+ bl_0_48 br_0_48 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c48
*+ bl_0_48 br_0_48 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c48
*+ bl_0_48 br_0_48 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c48
*+ bl_0_48 br_0_48 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c48
*+ bl_0_48 br_0_48 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c48
*+ bl_0_48 br_0_48 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c48
*+ bl_0_48 br_0_48 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c48
*+ bl_0_48 br_0_48 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c48
*+ bl_0_48 br_0_48 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c48
*+ bl_0_48 br_0_48 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c48
*+ bl_0_48 br_0_48 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c48
*+ bl_0_48 br_0_48 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c48
*+ bl_0_48 br_0_48 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c48
*+ bl_0_48 br_0_48 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c48
*+ bl_0_48 br_0_48 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c48
*+ bl_0_48 br_0_48 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c48
*+ bl_0_48 br_0_48 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c48
*+ bl_0_48 br_0_48 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c48
*+ bl_0_48 br_0_48 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c48
*+ bl_0_48 br_0_48 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c48
*+ bl_0_48 br_0_48 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c48
*+ bl_0_48 br_0_48 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c48
*+ bl_0_48 br_0_48 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c48
*+ bl_0_48 br_0_48 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c48
*+ bl_0_48 br_0_48 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c48
*+ bl_0_48 br_0_48 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c48
+ bl_0_48 br_0_48 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c49
+ bl_0_49 br_0_49 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c49
*+ bl_0_49 br_0_49 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c49
*+ bl_0_49 br_0_49 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c49
*+ bl_0_49 br_0_49 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c49
*+ bl_0_49 br_0_49 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c49
*+ bl_0_49 br_0_49 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c49
*+ bl_0_49 br_0_49 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c49
*+ bl_0_49 br_0_49 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c49
*+ bl_0_49 br_0_49 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c49
*+ bl_0_49 br_0_49 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c49
*+ bl_0_49 br_0_49 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c49
*+ bl_0_49 br_0_49 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c49
*+ bl_0_49 br_0_49 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c49
*+ bl_0_49 br_0_49 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c49
*+ bl_0_49 br_0_49 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c49
*+ bl_0_49 br_0_49 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c49
*+ bl_0_49 br_0_49 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c49
*+ bl_0_49 br_0_49 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c49
*+ bl_0_49 br_0_49 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c49
*+ bl_0_49 br_0_49 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c49
*+ bl_0_49 br_0_49 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c49
*+ bl_0_49 br_0_49 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c49
*+ bl_0_49 br_0_49 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c49
*+ bl_0_49 br_0_49 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c49
*+ bl_0_49 br_0_49 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c49
*+ bl_0_49 br_0_49 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c49
*+ bl_0_49 br_0_49 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c49
*+ bl_0_49 br_0_49 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c49
*+ bl_0_49 br_0_49 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c49
*+ bl_0_49 br_0_49 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c49
*+ bl_0_49 br_0_49 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c49
*+ bl_0_49 br_0_49 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c49
*+ bl_0_49 br_0_49 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c49
*+ bl_0_49 br_0_49 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c49
*+ bl_0_49 br_0_49 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c49
*+ bl_0_49 br_0_49 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c49
*+ bl_0_49 br_0_49 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c49
*+ bl_0_49 br_0_49 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c49
*+ bl_0_49 br_0_49 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c49
*+ bl_0_49 br_0_49 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c49
*+ bl_0_49 br_0_49 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c49
*+ bl_0_49 br_0_49 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c49
*+ bl_0_49 br_0_49 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c49
*+ bl_0_49 br_0_49 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c49
*+ bl_0_49 br_0_49 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c49
*+ bl_0_49 br_0_49 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c49
*+ bl_0_49 br_0_49 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c49
*+ bl_0_49 br_0_49 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c49
*+ bl_0_49 br_0_49 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c49
*+ bl_0_49 br_0_49 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c49
*+ bl_0_49 br_0_49 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c49
*+ bl_0_49 br_0_49 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c49
*+ bl_0_49 br_0_49 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c49
*+ bl_0_49 br_0_49 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c49
*+ bl_0_49 br_0_49 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c49
*+ bl_0_49 br_0_49 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c49
*+ bl_0_49 br_0_49 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c49
*+ bl_0_49 br_0_49 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c49
*+ bl_0_49 br_0_49 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c49
*+ bl_0_49 br_0_49 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c49
*+ bl_0_49 br_0_49 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c49
*+ bl_0_49 br_0_49 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c49
*+ bl_0_49 br_0_49 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c49
*+ bl_0_49 br_0_49 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c49
*+ bl_0_49 br_0_49 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c49
*+ bl_0_49 br_0_49 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c49
*+ bl_0_49 br_0_49 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c49
*+ bl_0_49 br_0_49 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c49
*+ bl_0_49 br_0_49 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c49
*+ bl_0_49 br_0_49 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c49
*+ bl_0_49 br_0_49 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c49
*+ bl_0_49 br_0_49 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c49
*+ bl_0_49 br_0_49 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c49
*+ bl_0_49 br_0_49 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c49
*+ bl_0_49 br_0_49 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c49
*+ bl_0_49 br_0_49 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c49
*+ bl_0_49 br_0_49 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c49
*+ bl_0_49 br_0_49 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c49
*+ bl_0_49 br_0_49 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c49
*+ bl_0_49 br_0_49 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c49
*+ bl_0_49 br_0_49 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c49
*+ bl_0_49 br_0_49 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c49
*+ bl_0_49 br_0_49 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c49
*+ bl_0_49 br_0_49 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c49
*+ bl_0_49 br_0_49 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c49
*+ bl_0_49 br_0_49 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c49
*+ bl_0_49 br_0_49 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c49
*+ bl_0_49 br_0_49 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c49
*+ bl_0_49 br_0_49 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c49
*+ bl_0_49 br_0_49 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c49
*+ bl_0_49 br_0_49 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c49
*+ bl_0_49 br_0_49 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c49
*+ bl_0_49 br_0_49 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c49
*+ bl_0_49 br_0_49 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c49
*+ bl_0_49 br_0_49 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c49
*+ bl_0_49 br_0_49 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c49
*+ bl_0_49 br_0_49 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c49
*+ bl_0_49 br_0_49 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c49
*+ bl_0_49 br_0_49 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c49
*+ bl_0_49 br_0_49 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c49
*+ bl_0_49 br_0_49 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c49
*+ bl_0_49 br_0_49 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c49
*+ bl_0_49 br_0_49 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c49
*+ bl_0_49 br_0_49 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c49
*+ bl_0_49 br_0_49 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c49
*+ bl_0_49 br_0_49 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c49
*+ bl_0_49 br_0_49 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c49
*+ bl_0_49 br_0_49 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c49
*+ bl_0_49 br_0_49 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c49
*+ bl_0_49 br_0_49 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c49
*+ bl_0_49 br_0_49 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c49
*+ bl_0_49 br_0_49 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c49
*+ bl_0_49 br_0_49 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c49
*+ bl_0_49 br_0_49 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c49
*+ bl_0_49 br_0_49 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c49
*+ bl_0_49 br_0_49 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c49
*+ bl_0_49 br_0_49 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c49
*+ bl_0_49 br_0_49 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c49
*+ bl_0_49 br_0_49 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c49
*+ bl_0_49 br_0_49 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c49
*+ bl_0_49 br_0_49 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c49
*+ bl_0_49 br_0_49 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c49
*+ bl_0_49 br_0_49 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c49
*+ bl_0_49 br_0_49 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c49
*+ bl_0_49 br_0_49 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c49
*+ bl_0_49 br_0_49 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c49
*+ bl_0_49 br_0_49 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c49
+ bl_0_49 br_0_49 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c50
+ bl_0_50 br_0_50 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c50
*+ bl_0_50 br_0_50 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c50
*+ bl_0_50 br_0_50 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c50
*+ bl_0_50 br_0_50 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c50
*+ bl_0_50 br_0_50 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c50
*+ bl_0_50 br_0_50 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c50
*+ bl_0_50 br_0_50 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c50
*+ bl_0_50 br_0_50 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c50
*+ bl_0_50 br_0_50 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c50
*+ bl_0_50 br_0_50 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c50
*+ bl_0_50 br_0_50 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c50
*+ bl_0_50 br_0_50 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c50
*+ bl_0_50 br_0_50 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c50
*+ bl_0_50 br_0_50 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c50
*+ bl_0_50 br_0_50 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c50
*+ bl_0_50 br_0_50 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c50
*+ bl_0_50 br_0_50 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c50
*+ bl_0_50 br_0_50 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c50
*+ bl_0_50 br_0_50 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c50
*+ bl_0_50 br_0_50 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c50
*+ bl_0_50 br_0_50 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c50
*+ bl_0_50 br_0_50 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c50
*+ bl_0_50 br_0_50 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c50
*+ bl_0_50 br_0_50 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c50
*+ bl_0_50 br_0_50 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c50
*+ bl_0_50 br_0_50 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c50
*+ bl_0_50 br_0_50 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c50
*+ bl_0_50 br_0_50 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c50
*+ bl_0_50 br_0_50 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c50
*+ bl_0_50 br_0_50 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c50
*+ bl_0_50 br_0_50 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c50
*+ bl_0_50 br_0_50 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c50
*+ bl_0_50 br_0_50 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c50
*+ bl_0_50 br_0_50 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c50
*+ bl_0_50 br_0_50 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c50
*+ bl_0_50 br_0_50 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c50
*+ bl_0_50 br_0_50 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c50
*+ bl_0_50 br_0_50 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c50
*+ bl_0_50 br_0_50 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c50
*+ bl_0_50 br_0_50 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c50
*+ bl_0_50 br_0_50 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c50
*+ bl_0_50 br_0_50 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c50
*+ bl_0_50 br_0_50 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c50
*+ bl_0_50 br_0_50 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c50
*+ bl_0_50 br_0_50 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c50
*+ bl_0_50 br_0_50 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c50
*+ bl_0_50 br_0_50 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c50
*+ bl_0_50 br_0_50 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c50
*+ bl_0_50 br_0_50 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c50
*+ bl_0_50 br_0_50 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c50
*+ bl_0_50 br_0_50 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c50
*+ bl_0_50 br_0_50 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c50
*+ bl_0_50 br_0_50 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c50
*+ bl_0_50 br_0_50 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c50
*+ bl_0_50 br_0_50 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c50
*+ bl_0_50 br_0_50 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c50
*+ bl_0_50 br_0_50 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c50
*+ bl_0_50 br_0_50 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c50
*+ bl_0_50 br_0_50 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c50
*+ bl_0_50 br_0_50 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c50
*+ bl_0_50 br_0_50 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c50
*+ bl_0_50 br_0_50 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c50
*+ bl_0_50 br_0_50 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c50
*+ bl_0_50 br_0_50 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c50
*+ bl_0_50 br_0_50 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c50
*+ bl_0_50 br_0_50 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c50
*+ bl_0_50 br_0_50 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c50
*+ bl_0_50 br_0_50 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c50
*+ bl_0_50 br_0_50 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c50
*+ bl_0_50 br_0_50 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c50
*+ bl_0_50 br_0_50 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c50
*+ bl_0_50 br_0_50 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c50
*+ bl_0_50 br_0_50 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c50
*+ bl_0_50 br_0_50 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c50
*+ bl_0_50 br_0_50 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c50
*+ bl_0_50 br_0_50 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c50
*+ bl_0_50 br_0_50 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c50
*+ bl_0_50 br_0_50 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c50
*+ bl_0_50 br_0_50 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c50
*+ bl_0_50 br_0_50 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c50
*+ bl_0_50 br_0_50 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c50
*+ bl_0_50 br_0_50 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c50
*+ bl_0_50 br_0_50 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c50
*+ bl_0_50 br_0_50 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c50
*+ bl_0_50 br_0_50 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c50
*+ bl_0_50 br_0_50 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c50
*+ bl_0_50 br_0_50 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c50
*+ bl_0_50 br_0_50 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c50
*+ bl_0_50 br_0_50 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c50
*+ bl_0_50 br_0_50 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c50
*+ bl_0_50 br_0_50 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c50
*+ bl_0_50 br_0_50 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c50
*+ bl_0_50 br_0_50 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c50
*+ bl_0_50 br_0_50 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c50
*+ bl_0_50 br_0_50 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c50
*+ bl_0_50 br_0_50 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c50
*+ bl_0_50 br_0_50 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c50
*+ bl_0_50 br_0_50 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c50
*+ bl_0_50 br_0_50 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c50
*+ bl_0_50 br_0_50 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c50
*+ bl_0_50 br_0_50 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c50
*+ bl_0_50 br_0_50 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c50
*+ bl_0_50 br_0_50 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c50
*+ bl_0_50 br_0_50 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c50
*+ bl_0_50 br_0_50 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c50
*+ bl_0_50 br_0_50 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c50
*+ bl_0_50 br_0_50 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c50
*+ bl_0_50 br_0_50 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c50
*+ bl_0_50 br_0_50 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c50
*+ bl_0_50 br_0_50 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c50
*+ bl_0_50 br_0_50 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c50
*+ bl_0_50 br_0_50 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c50
*+ bl_0_50 br_0_50 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c50
*+ bl_0_50 br_0_50 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c50
*+ bl_0_50 br_0_50 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c50
*+ bl_0_50 br_0_50 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c50
*+ bl_0_50 br_0_50 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c50
*+ bl_0_50 br_0_50 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c50
*+ bl_0_50 br_0_50 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c50
*+ bl_0_50 br_0_50 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c50
*+ bl_0_50 br_0_50 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c50
*+ bl_0_50 br_0_50 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c50
*+ bl_0_50 br_0_50 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c50
*+ bl_0_50 br_0_50 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c50
*+ bl_0_50 br_0_50 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c50
*+ bl_0_50 br_0_50 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c50
*+ bl_0_50 br_0_50 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c50
+ bl_0_50 br_0_50 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c51
+ bl_0_51 br_0_51 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c51
*+ bl_0_51 br_0_51 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c51
*+ bl_0_51 br_0_51 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c51
*+ bl_0_51 br_0_51 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c51
*+ bl_0_51 br_0_51 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c51
*+ bl_0_51 br_0_51 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c51
*+ bl_0_51 br_0_51 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c51
*+ bl_0_51 br_0_51 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c51
*+ bl_0_51 br_0_51 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c51
*+ bl_0_51 br_0_51 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c51
*+ bl_0_51 br_0_51 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c51
*+ bl_0_51 br_0_51 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c51
*+ bl_0_51 br_0_51 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c51
*+ bl_0_51 br_0_51 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c51
*+ bl_0_51 br_0_51 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c51
*+ bl_0_51 br_0_51 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c51
*+ bl_0_51 br_0_51 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c51
*+ bl_0_51 br_0_51 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c51
*+ bl_0_51 br_0_51 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c51
*+ bl_0_51 br_0_51 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c51
*+ bl_0_51 br_0_51 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c51
*+ bl_0_51 br_0_51 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c51
*+ bl_0_51 br_0_51 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c51
*+ bl_0_51 br_0_51 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c51
*+ bl_0_51 br_0_51 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c51
*+ bl_0_51 br_0_51 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c51
*+ bl_0_51 br_0_51 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c51
*+ bl_0_51 br_0_51 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c51
*+ bl_0_51 br_0_51 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c51
*+ bl_0_51 br_0_51 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c51
*+ bl_0_51 br_0_51 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c51
*+ bl_0_51 br_0_51 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c51
*+ bl_0_51 br_0_51 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c51
*+ bl_0_51 br_0_51 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c51
*+ bl_0_51 br_0_51 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c51
*+ bl_0_51 br_0_51 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c51
*+ bl_0_51 br_0_51 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c51
*+ bl_0_51 br_0_51 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c51
*+ bl_0_51 br_0_51 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c51
*+ bl_0_51 br_0_51 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c51
*+ bl_0_51 br_0_51 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c51
*+ bl_0_51 br_0_51 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c51
*+ bl_0_51 br_0_51 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c51
*+ bl_0_51 br_0_51 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c51
*+ bl_0_51 br_0_51 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c51
*+ bl_0_51 br_0_51 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c51
*+ bl_0_51 br_0_51 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c51
*+ bl_0_51 br_0_51 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c51
*+ bl_0_51 br_0_51 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c51
*+ bl_0_51 br_0_51 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c51
*+ bl_0_51 br_0_51 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c51
*+ bl_0_51 br_0_51 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c51
*+ bl_0_51 br_0_51 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c51
*+ bl_0_51 br_0_51 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c51
*+ bl_0_51 br_0_51 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c51
*+ bl_0_51 br_0_51 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c51
*+ bl_0_51 br_0_51 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c51
*+ bl_0_51 br_0_51 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c51
*+ bl_0_51 br_0_51 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c51
*+ bl_0_51 br_0_51 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c51
*+ bl_0_51 br_0_51 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c51
*+ bl_0_51 br_0_51 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c51
*+ bl_0_51 br_0_51 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c51
*+ bl_0_51 br_0_51 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c51
*+ bl_0_51 br_0_51 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c51
*+ bl_0_51 br_0_51 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c51
*+ bl_0_51 br_0_51 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c51
*+ bl_0_51 br_0_51 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c51
*+ bl_0_51 br_0_51 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c51
*+ bl_0_51 br_0_51 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c51
*+ bl_0_51 br_0_51 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c51
*+ bl_0_51 br_0_51 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c51
*+ bl_0_51 br_0_51 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c51
*+ bl_0_51 br_0_51 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c51
*+ bl_0_51 br_0_51 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c51
*+ bl_0_51 br_0_51 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c51
*+ bl_0_51 br_0_51 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c51
*+ bl_0_51 br_0_51 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c51
*+ bl_0_51 br_0_51 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c51
*+ bl_0_51 br_0_51 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c51
*+ bl_0_51 br_0_51 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c51
*+ bl_0_51 br_0_51 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c51
*+ bl_0_51 br_0_51 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c51
*+ bl_0_51 br_0_51 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c51
*+ bl_0_51 br_0_51 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c51
*+ bl_0_51 br_0_51 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c51
*+ bl_0_51 br_0_51 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c51
*+ bl_0_51 br_0_51 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c51
*+ bl_0_51 br_0_51 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c51
*+ bl_0_51 br_0_51 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c51
*+ bl_0_51 br_0_51 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c51
*+ bl_0_51 br_0_51 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c51
*+ bl_0_51 br_0_51 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c51
*+ bl_0_51 br_0_51 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c51
*+ bl_0_51 br_0_51 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c51
*+ bl_0_51 br_0_51 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c51
*+ bl_0_51 br_0_51 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c51
*+ bl_0_51 br_0_51 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c51
*+ bl_0_51 br_0_51 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c51
*+ bl_0_51 br_0_51 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c51
*+ bl_0_51 br_0_51 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c51
*+ bl_0_51 br_0_51 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c51
*+ bl_0_51 br_0_51 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c51
*+ bl_0_51 br_0_51 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c51
*+ bl_0_51 br_0_51 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c51
*+ bl_0_51 br_0_51 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c51
*+ bl_0_51 br_0_51 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c51
*+ bl_0_51 br_0_51 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c51
*+ bl_0_51 br_0_51 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c51
*+ bl_0_51 br_0_51 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c51
*+ bl_0_51 br_0_51 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c51
*+ bl_0_51 br_0_51 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c51
*+ bl_0_51 br_0_51 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c51
*+ bl_0_51 br_0_51 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c51
*+ bl_0_51 br_0_51 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c51
*+ bl_0_51 br_0_51 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c51
*+ bl_0_51 br_0_51 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c51
*+ bl_0_51 br_0_51 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c51
*+ bl_0_51 br_0_51 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c51
*+ bl_0_51 br_0_51 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c51
*+ bl_0_51 br_0_51 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c51
*+ bl_0_51 br_0_51 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c51
*+ bl_0_51 br_0_51 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c51
*+ bl_0_51 br_0_51 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c51
*+ bl_0_51 br_0_51 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c51
*+ bl_0_51 br_0_51 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c51
*+ bl_0_51 br_0_51 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c51
+ bl_0_51 br_0_51 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c52
+ bl_0_52 br_0_52 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c52
*+ bl_0_52 br_0_52 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c52
*+ bl_0_52 br_0_52 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c52
*+ bl_0_52 br_0_52 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c52
*+ bl_0_52 br_0_52 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c52
*+ bl_0_52 br_0_52 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c52
*+ bl_0_52 br_0_52 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c52
*+ bl_0_52 br_0_52 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c52
*+ bl_0_52 br_0_52 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c52
*+ bl_0_52 br_0_52 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c52
*+ bl_0_52 br_0_52 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c52
*+ bl_0_52 br_0_52 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c52
*+ bl_0_52 br_0_52 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c52
*+ bl_0_52 br_0_52 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c52
*+ bl_0_52 br_0_52 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c52
*+ bl_0_52 br_0_52 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c52
*+ bl_0_52 br_0_52 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c52
*+ bl_0_52 br_0_52 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c52
*+ bl_0_52 br_0_52 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c52
*+ bl_0_52 br_0_52 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c52
*+ bl_0_52 br_0_52 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c52
*+ bl_0_52 br_0_52 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c52
*+ bl_0_52 br_0_52 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c52
*+ bl_0_52 br_0_52 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c52
*+ bl_0_52 br_0_52 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c52
*+ bl_0_52 br_0_52 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c52
*+ bl_0_52 br_0_52 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c52
*+ bl_0_52 br_0_52 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c52
*+ bl_0_52 br_0_52 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c52
*+ bl_0_52 br_0_52 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c52
*+ bl_0_52 br_0_52 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c52
*+ bl_0_52 br_0_52 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c52
*+ bl_0_52 br_0_52 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c52
*+ bl_0_52 br_0_52 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c52
*+ bl_0_52 br_0_52 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c52
*+ bl_0_52 br_0_52 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c52
*+ bl_0_52 br_0_52 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c52
*+ bl_0_52 br_0_52 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c52
*+ bl_0_52 br_0_52 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c52
*+ bl_0_52 br_0_52 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c52
*+ bl_0_52 br_0_52 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c52
*+ bl_0_52 br_0_52 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c52
*+ bl_0_52 br_0_52 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c52
*+ bl_0_52 br_0_52 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c52
*+ bl_0_52 br_0_52 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c52
*+ bl_0_52 br_0_52 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c52
*+ bl_0_52 br_0_52 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c52
*+ bl_0_52 br_0_52 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c52
*+ bl_0_52 br_0_52 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c52
*+ bl_0_52 br_0_52 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c52
*+ bl_0_52 br_0_52 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c52
*+ bl_0_52 br_0_52 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c52
*+ bl_0_52 br_0_52 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c52
*+ bl_0_52 br_0_52 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c52
*+ bl_0_52 br_0_52 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c52
*+ bl_0_52 br_0_52 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c52
*+ bl_0_52 br_0_52 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c52
*+ bl_0_52 br_0_52 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c52
*+ bl_0_52 br_0_52 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c52
*+ bl_0_52 br_0_52 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c52
*+ bl_0_52 br_0_52 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c52
*+ bl_0_52 br_0_52 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c52
*+ bl_0_52 br_0_52 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c52
*+ bl_0_52 br_0_52 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c52
*+ bl_0_52 br_0_52 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c52
*+ bl_0_52 br_0_52 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c52
*+ bl_0_52 br_0_52 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c52
*+ bl_0_52 br_0_52 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c52
*+ bl_0_52 br_0_52 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c52
*+ bl_0_52 br_0_52 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c52
*+ bl_0_52 br_0_52 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c52
*+ bl_0_52 br_0_52 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c52
*+ bl_0_52 br_0_52 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c52
*+ bl_0_52 br_0_52 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c52
*+ bl_0_52 br_0_52 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c52
*+ bl_0_52 br_0_52 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c52
*+ bl_0_52 br_0_52 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c52
*+ bl_0_52 br_0_52 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c52
*+ bl_0_52 br_0_52 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c52
*+ bl_0_52 br_0_52 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c52
*+ bl_0_52 br_0_52 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c52
*+ bl_0_52 br_0_52 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c52
*+ bl_0_52 br_0_52 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c52
*+ bl_0_52 br_0_52 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c52
*+ bl_0_52 br_0_52 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c52
*+ bl_0_52 br_0_52 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c52
*+ bl_0_52 br_0_52 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c52
*+ bl_0_52 br_0_52 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c52
*+ bl_0_52 br_0_52 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c52
*+ bl_0_52 br_0_52 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c52
*+ bl_0_52 br_0_52 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c52
*+ bl_0_52 br_0_52 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c52
*+ bl_0_52 br_0_52 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c52
*+ bl_0_52 br_0_52 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c52
*+ bl_0_52 br_0_52 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c52
*+ bl_0_52 br_0_52 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c52
*+ bl_0_52 br_0_52 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c52
*+ bl_0_52 br_0_52 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c52
*+ bl_0_52 br_0_52 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c52
*+ bl_0_52 br_0_52 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c52
*+ bl_0_52 br_0_52 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c52
*+ bl_0_52 br_0_52 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c52
*+ bl_0_52 br_0_52 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c52
*+ bl_0_52 br_0_52 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c52
*+ bl_0_52 br_0_52 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c52
*+ bl_0_52 br_0_52 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c52
*+ bl_0_52 br_0_52 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c52
*+ bl_0_52 br_0_52 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c52
*+ bl_0_52 br_0_52 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c52
*+ bl_0_52 br_0_52 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c52
*+ bl_0_52 br_0_52 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c52
*+ bl_0_52 br_0_52 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c52
*+ bl_0_52 br_0_52 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c52
*+ bl_0_52 br_0_52 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c52
*+ bl_0_52 br_0_52 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c52
*+ bl_0_52 br_0_52 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c52
*+ bl_0_52 br_0_52 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c52
*+ bl_0_52 br_0_52 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c52
*+ bl_0_52 br_0_52 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c52
*+ bl_0_52 br_0_52 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c52
*+ bl_0_52 br_0_52 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c52
*+ bl_0_52 br_0_52 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c52
*+ bl_0_52 br_0_52 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c52
*+ bl_0_52 br_0_52 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c52
*+ bl_0_52 br_0_52 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c52
*+ bl_0_52 br_0_52 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c52
*+ bl_0_52 br_0_52 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c52
+ bl_0_52 br_0_52 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c53
+ bl_0_53 br_0_53 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c53
*+ bl_0_53 br_0_53 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c53
*+ bl_0_53 br_0_53 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c53
*+ bl_0_53 br_0_53 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c53
*+ bl_0_53 br_0_53 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c53
*+ bl_0_53 br_0_53 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c53
*+ bl_0_53 br_0_53 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c53
*+ bl_0_53 br_0_53 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c53
*+ bl_0_53 br_0_53 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c53
*+ bl_0_53 br_0_53 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c53
*+ bl_0_53 br_0_53 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c53
*+ bl_0_53 br_0_53 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c53
*+ bl_0_53 br_0_53 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c53
*+ bl_0_53 br_0_53 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c53
*+ bl_0_53 br_0_53 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c53
*+ bl_0_53 br_0_53 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c53
*+ bl_0_53 br_0_53 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c53
*+ bl_0_53 br_0_53 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c53
*+ bl_0_53 br_0_53 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c53
*+ bl_0_53 br_0_53 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c53
*+ bl_0_53 br_0_53 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c53
*+ bl_0_53 br_0_53 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c53
*+ bl_0_53 br_0_53 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c53
*+ bl_0_53 br_0_53 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c53
*+ bl_0_53 br_0_53 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c53
*+ bl_0_53 br_0_53 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c53
*+ bl_0_53 br_0_53 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c53
*+ bl_0_53 br_0_53 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c53
*+ bl_0_53 br_0_53 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c53
*+ bl_0_53 br_0_53 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c53
*+ bl_0_53 br_0_53 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c53
*+ bl_0_53 br_0_53 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c53
*+ bl_0_53 br_0_53 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c53
*+ bl_0_53 br_0_53 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c53
*+ bl_0_53 br_0_53 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c53
*+ bl_0_53 br_0_53 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c53
*+ bl_0_53 br_0_53 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c53
*+ bl_0_53 br_0_53 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c53
*+ bl_0_53 br_0_53 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c53
*+ bl_0_53 br_0_53 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c53
*+ bl_0_53 br_0_53 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c53
*+ bl_0_53 br_0_53 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c53
*+ bl_0_53 br_0_53 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c53
*+ bl_0_53 br_0_53 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c53
*+ bl_0_53 br_0_53 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c53
*+ bl_0_53 br_0_53 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c53
*+ bl_0_53 br_0_53 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c53
*+ bl_0_53 br_0_53 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c53
*+ bl_0_53 br_0_53 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c53
*+ bl_0_53 br_0_53 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c53
*+ bl_0_53 br_0_53 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c53
*+ bl_0_53 br_0_53 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c53
*+ bl_0_53 br_0_53 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c53
*+ bl_0_53 br_0_53 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c53
*+ bl_0_53 br_0_53 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c53
*+ bl_0_53 br_0_53 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c53
*+ bl_0_53 br_0_53 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c53
*+ bl_0_53 br_0_53 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c53
*+ bl_0_53 br_0_53 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c53
*+ bl_0_53 br_0_53 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c53
*+ bl_0_53 br_0_53 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c53
*+ bl_0_53 br_0_53 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c53
*+ bl_0_53 br_0_53 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c53
*+ bl_0_53 br_0_53 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c53
*+ bl_0_53 br_0_53 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c53
*+ bl_0_53 br_0_53 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c53
*+ bl_0_53 br_0_53 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c53
*+ bl_0_53 br_0_53 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c53
*+ bl_0_53 br_0_53 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c53
*+ bl_0_53 br_0_53 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c53
*+ bl_0_53 br_0_53 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c53
*+ bl_0_53 br_0_53 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c53
*+ bl_0_53 br_0_53 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c53
*+ bl_0_53 br_0_53 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c53
*+ bl_0_53 br_0_53 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c53
*+ bl_0_53 br_0_53 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c53
*+ bl_0_53 br_0_53 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c53
*+ bl_0_53 br_0_53 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c53
*+ bl_0_53 br_0_53 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c53
*+ bl_0_53 br_0_53 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c53
*+ bl_0_53 br_0_53 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c53
*+ bl_0_53 br_0_53 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c53
*+ bl_0_53 br_0_53 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c53
*+ bl_0_53 br_0_53 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c53
*+ bl_0_53 br_0_53 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c53
*+ bl_0_53 br_0_53 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c53
*+ bl_0_53 br_0_53 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c53
*+ bl_0_53 br_0_53 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c53
*+ bl_0_53 br_0_53 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c53
*+ bl_0_53 br_0_53 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c53
*+ bl_0_53 br_0_53 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c53
*+ bl_0_53 br_0_53 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c53
*+ bl_0_53 br_0_53 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c53
*+ bl_0_53 br_0_53 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c53
*+ bl_0_53 br_0_53 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c53
*+ bl_0_53 br_0_53 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c53
*+ bl_0_53 br_0_53 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c53
*+ bl_0_53 br_0_53 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c53
*+ bl_0_53 br_0_53 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c53
*+ bl_0_53 br_0_53 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c53
*+ bl_0_53 br_0_53 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c53
*+ bl_0_53 br_0_53 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c53
*+ bl_0_53 br_0_53 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c53
*+ bl_0_53 br_0_53 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c53
*+ bl_0_53 br_0_53 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c53
*+ bl_0_53 br_0_53 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c53
*+ bl_0_53 br_0_53 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c53
*+ bl_0_53 br_0_53 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c53
*+ bl_0_53 br_0_53 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c53
*+ bl_0_53 br_0_53 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c53
*+ bl_0_53 br_0_53 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c53
*+ bl_0_53 br_0_53 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c53
*+ bl_0_53 br_0_53 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c53
*+ bl_0_53 br_0_53 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c53
*+ bl_0_53 br_0_53 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c53
*+ bl_0_53 br_0_53 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c53
*+ bl_0_53 br_0_53 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c53
*+ bl_0_53 br_0_53 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c53
*+ bl_0_53 br_0_53 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c53
*+ bl_0_53 br_0_53 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c53
*+ bl_0_53 br_0_53 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c53
*+ bl_0_53 br_0_53 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c53
*+ bl_0_53 br_0_53 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c53
*+ bl_0_53 br_0_53 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c53
*+ bl_0_53 br_0_53 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c53
*+ bl_0_53 br_0_53 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c53
*+ bl_0_53 br_0_53 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c53
+ bl_0_53 br_0_53 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c54
+ bl_0_54 br_0_54 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c54
*+ bl_0_54 br_0_54 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c54
*+ bl_0_54 br_0_54 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c54
*+ bl_0_54 br_0_54 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c54
*+ bl_0_54 br_0_54 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c54
*+ bl_0_54 br_0_54 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c54
*+ bl_0_54 br_0_54 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c54
*+ bl_0_54 br_0_54 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c54
*+ bl_0_54 br_0_54 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c54
*+ bl_0_54 br_0_54 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c54
*+ bl_0_54 br_0_54 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c54
*+ bl_0_54 br_0_54 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c54
*+ bl_0_54 br_0_54 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c54
*+ bl_0_54 br_0_54 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c54
*+ bl_0_54 br_0_54 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c54
*+ bl_0_54 br_0_54 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c54
*+ bl_0_54 br_0_54 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c54
*+ bl_0_54 br_0_54 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c54
*+ bl_0_54 br_0_54 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c54
*+ bl_0_54 br_0_54 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c54
*+ bl_0_54 br_0_54 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c54
*+ bl_0_54 br_0_54 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c54
*+ bl_0_54 br_0_54 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c54
*+ bl_0_54 br_0_54 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c54
*+ bl_0_54 br_0_54 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c54
*+ bl_0_54 br_0_54 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c54
*+ bl_0_54 br_0_54 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c54
*+ bl_0_54 br_0_54 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c54
*+ bl_0_54 br_0_54 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c54
*+ bl_0_54 br_0_54 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c54
*+ bl_0_54 br_0_54 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c54
*+ bl_0_54 br_0_54 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c54
*+ bl_0_54 br_0_54 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c54
*+ bl_0_54 br_0_54 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c54
*+ bl_0_54 br_0_54 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c54
*+ bl_0_54 br_0_54 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c54
*+ bl_0_54 br_0_54 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c54
*+ bl_0_54 br_0_54 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c54
*+ bl_0_54 br_0_54 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c54
*+ bl_0_54 br_0_54 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c54
*+ bl_0_54 br_0_54 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c54
*+ bl_0_54 br_0_54 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c54
*+ bl_0_54 br_0_54 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c54
*+ bl_0_54 br_0_54 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c54
*+ bl_0_54 br_0_54 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c54
*+ bl_0_54 br_0_54 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c54
*+ bl_0_54 br_0_54 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c54
*+ bl_0_54 br_0_54 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c54
*+ bl_0_54 br_0_54 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c54
*+ bl_0_54 br_0_54 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c54
*+ bl_0_54 br_0_54 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c54
*+ bl_0_54 br_0_54 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c54
*+ bl_0_54 br_0_54 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c54
*+ bl_0_54 br_0_54 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c54
*+ bl_0_54 br_0_54 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c54
*+ bl_0_54 br_0_54 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c54
*+ bl_0_54 br_0_54 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c54
*+ bl_0_54 br_0_54 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c54
*+ bl_0_54 br_0_54 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c54
*+ bl_0_54 br_0_54 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c54
*+ bl_0_54 br_0_54 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c54
*+ bl_0_54 br_0_54 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c54
*+ bl_0_54 br_0_54 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c54
*+ bl_0_54 br_0_54 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c54
*+ bl_0_54 br_0_54 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c54
*+ bl_0_54 br_0_54 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c54
*+ bl_0_54 br_0_54 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c54
*+ bl_0_54 br_0_54 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c54
*+ bl_0_54 br_0_54 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c54
*+ bl_0_54 br_0_54 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c54
*+ bl_0_54 br_0_54 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c54
*+ bl_0_54 br_0_54 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c54
*+ bl_0_54 br_0_54 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c54
*+ bl_0_54 br_0_54 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c54
*+ bl_0_54 br_0_54 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c54
*+ bl_0_54 br_0_54 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c54
*+ bl_0_54 br_0_54 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c54
*+ bl_0_54 br_0_54 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c54
*+ bl_0_54 br_0_54 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c54
*+ bl_0_54 br_0_54 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c54
*+ bl_0_54 br_0_54 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c54
*+ bl_0_54 br_0_54 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c54
*+ bl_0_54 br_0_54 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c54
*+ bl_0_54 br_0_54 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c54
*+ bl_0_54 br_0_54 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c54
*+ bl_0_54 br_0_54 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c54
*+ bl_0_54 br_0_54 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c54
*+ bl_0_54 br_0_54 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c54
*+ bl_0_54 br_0_54 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c54
*+ bl_0_54 br_0_54 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c54
*+ bl_0_54 br_0_54 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c54
*+ bl_0_54 br_0_54 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c54
*+ bl_0_54 br_0_54 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c54
*+ bl_0_54 br_0_54 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c54
*+ bl_0_54 br_0_54 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c54
*+ bl_0_54 br_0_54 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c54
*+ bl_0_54 br_0_54 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c54
*+ bl_0_54 br_0_54 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c54
*+ bl_0_54 br_0_54 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c54
*+ bl_0_54 br_0_54 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c54
*+ bl_0_54 br_0_54 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c54
*+ bl_0_54 br_0_54 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c54
*+ bl_0_54 br_0_54 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c54
*+ bl_0_54 br_0_54 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c54
*+ bl_0_54 br_0_54 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c54
*+ bl_0_54 br_0_54 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c54
*+ bl_0_54 br_0_54 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c54
*+ bl_0_54 br_0_54 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c54
*+ bl_0_54 br_0_54 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c54
*+ bl_0_54 br_0_54 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c54
*+ bl_0_54 br_0_54 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c54
*+ bl_0_54 br_0_54 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c54
*+ bl_0_54 br_0_54 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c54
*+ bl_0_54 br_0_54 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c54
*+ bl_0_54 br_0_54 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c54
*+ bl_0_54 br_0_54 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c54
*+ bl_0_54 br_0_54 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c54
*+ bl_0_54 br_0_54 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c54
*+ bl_0_54 br_0_54 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c54
*+ bl_0_54 br_0_54 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c54
*+ bl_0_54 br_0_54 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c54
*+ bl_0_54 br_0_54 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c54
*+ bl_0_54 br_0_54 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c54
*+ bl_0_54 br_0_54 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c54
*+ bl_0_54 br_0_54 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c54
*+ bl_0_54 br_0_54 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c54
*+ bl_0_54 br_0_54 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c54
+ bl_0_54 br_0_54 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c55
+ bl_0_55 br_0_55 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c55
*+ bl_0_55 br_0_55 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c55
*+ bl_0_55 br_0_55 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c55
*+ bl_0_55 br_0_55 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c55
*+ bl_0_55 br_0_55 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c55
*+ bl_0_55 br_0_55 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c55
*+ bl_0_55 br_0_55 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c55
*+ bl_0_55 br_0_55 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c55
*+ bl_0_55 br_0_55 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c55
*+ bl_0_55 br_0_55 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c55
*+ bl_0_55 br_0_55 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c55
*+ bl_0_55 br_0_55 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c55
*+ bl_0_55 br_0_55 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c55
*+ bl_0_55 br_0_55 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c55
*+ bl_0_55 br_0_55 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c55
*+ bl_0_55 br_0_55 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c55
*+ bl_0_55 br_0_55 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c55
*+ bl_0_55 br_0_55 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c55
*+ bl_0_55 br_0_55 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c55
*+ bl_0_55 br_0_55 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c55
*+ bl_0_55 br_0_55 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c55
*+ bl_0_55 br_0_55 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c55
*+ bl_0_55 br_0_55 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c55
*+ bl_0_55 br_0_55 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c55
*+ bl_0_55 br_0_55 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c55
*+ bl_0_55 br_0_55 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c55
*+ bl_0_55 br_0_55 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c55
*+ bl_0_55 br_0_55 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c55
*+ bl_0_55 br_0_55 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c55
*+ bl_0_55 br_0_55 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c55
*+ bl_0_55 br_0_55 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c55
*+ bl_0_55 br_0_55 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c55
*+ bl_0_55 br_0_55 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c55
*+ bl_0_55 br_0_55 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c55
*+ bl_0_55 br_0_55 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c55
*+ bl_0_55 br_0_55 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c55
*+ bl_0_55 br_0_55 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c55
*+ bl_0_55 br_0_55 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c55
*+ bl_0_55 br_0_55 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c55
*+ bl_0_55 br_0_55 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c55
*+ bl_0_55 br_0_55 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c55
*+ bl_0_55 br_0_55 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c55
*+ bl_0_55 br_0_55 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c55
*+ bl_0_55 br_0_55 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c55
*+ bl_0_55 br_0_55 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c55
*+ bl_0_55 br_0_55 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c55
*+ bl_0_55 br_0_55 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c55
*+ bl_0_55 br_0_55 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c55
*+ bl_0_55 br_0_55 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c55
*+ bl_0_55 br_0_55 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c55
*+ bl_0_55 br_0_55 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c55
*+ bl_0_55 br_0_55 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c55
*+ bl_0_55 br_0_55 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c55
*+ bl_0_55 br_0_55 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c55
*+ bl_0_55 br_0_55 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c55
*+ bl_0_55 br_0_55 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c55
*+ bl_0_55 br_0_55 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c55
*+ bl_0_55 br_0_55 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c55
*+ bl_0_55 br_0_55 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c55
*+ bl_0_55 br_0_55 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c55
*+ bl_0_55 br_0_55 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c55
*+ bl_0_55 br_0_55 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c55
*+ bl_0_55 br_0_55 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c55
*+ bl_0_55 br_0_55 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c55
*+ bl_0_55 br_0_55 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c55
*+ bl_0_55 br_0_55 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c55
*+ bl_0_55 br_0_55 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c55
*+ bl_0_55 br_0_55 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c55
*+ bl_0_55 br_0_55 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c55
*+ bl_0_55 br_0_55 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c55
*+ bl_0_55 br_0_55 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c55
*+ bl_0_55 br_0_55 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c55
*+ bl_0_55 br_0_55 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c55
*+ bl_0_55 br_0_55 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c55
*+ bl_0_55 br_0_55 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c55
*+ bl_0_55 br_0_55 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c55
*+ bl_0_55 br_0_55 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c55
*+ bl_0_55 br_0_55 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c55
*+ bl_0_55 br_0_55 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c55
*+ bl_0_55 br_0_55 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c55
*+ bl_0_55 br_0_55 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c55
*+ bl_0_55 br_0_55 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c55
*+ bl_0_55 br_0_55 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c55
*+ bl_0_55 br_0_55 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c55
*+ bl_0_55 br_0_55 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c55
*+ bl_0_55 br_0_55 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c55
*+ bl_0_55 br_0_55 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c55
*+ bl_0_55 br_0_55 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c55
*+ bl_0_55 br_0_55 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c55
*+ bl_0_55 br_0_55 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c55
*+ bl_0_55 br_0_55 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c55
*+ bl_0_55 br_0_55 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c55
*+ bl_0_55 br_0_55 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c55
*+ bl_0_55 br_0_55 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c55
*+ bl_0_55 br_0_55 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c55
*+ bl_0_55 br_0_55 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c55
*+ bl_0_55 br_0_55 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c55
*+ bl_0_55 br_0_55 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c55
*+ bl_0_55 br_0_55 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c55
*+ bl_0_55 br_0_55 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c55
*+ bl_0_55 br_0_55 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c55
*+ bl_0_55 br_0_55 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c55
*+ bl_0_55 br_0_55 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c55
*+ bl_0_55 br_0_55 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c55
*+ bl_0_55 br_0_55 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c55
*+ bl_0_55 br_0_55 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c55
*+ bl_0_55 br_0_55 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c55
*+ bl_0_55 br_0_55 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c55
*+ bl_0_55 br_0_55 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c55
*+ bl_0_55 br_0_55 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c55
*+ bl_0_55 br_0_55 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c55
*+ bl_0_55 br_0_55 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c55
*+ bl_0_55 br_0_55 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c55
*+ bl_0_55 br_0_55 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c55
*+ bl_0_55 br_0_55 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c55
*+ bl_0_55 br_0_55 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c55
*+ bl_0_55 br_0_55 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c55
*+ bl_0_55 br_0_55 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c55
*+ bl_0_55 br_0_55 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c55
*+ bl_0_55 br_0_55 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c55
*+ bl_0_55 br_0_55 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c55
*+ bl_0_55 br_0_55 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c55
*+ bl_0_55 br_0_55 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c55
*+ bl_0_55 br_0_55 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c55
*+ bl_0_55 br_0_55 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c55
*+ bl_0_55 br_0_55 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c55
*+ bl_0_55 br_0_55 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c55
+ bl_0_55 br_0_55 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c56
+ bl_0_56 br_0_56 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c56
*+ bl_0_56 br_0_56 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c56
*+ bl_0_56 br_0_56 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c56
*+ bl_0_56 br_0_56 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c56
*+ bl_0_56 br_0_56 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c56
*+ bl_0_56 br_0_56 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c56
*+ bl_0_56 br_0_56 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c56
*+ bl_0_56 br_0_56 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c56
*+ bl_0_56 br_0_56 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c56
*+ bl_0_56 br_0_56 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c56
*+ bl_0_56 br_0_56 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c56
*+ bl_0_56 br_0_56 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c56
*+ bl_0_56 br_0_56 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c56
*+ bl_0_56 br_0_56 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c56
*+ bl_0_56 br_0_56 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c56
*+ bl_0_56 br_0_56 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c56
*+ bl_0_56 br_0_56 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c56
*+ bl_0_56 br_0_56 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c56
*+ bl_0_56 br_0_56 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c56
*+ bl_0_56 br_0_56 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c56
*+ bl_0_56 br_0_56 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c56
*+ bl_0_56 br_0_56 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c56
*+ bl_0_56 br_0_56 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c56
*+ bl_0_56 br_0_56 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c56
*+ bl_0_56 br_0_56 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c56
*+ bl_0_56 br_0_56 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c56
*+ bl_0_56 br_0_56 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c56
*+ bl_0_56 br_0_56 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c56
*+ bl_0_56 br_0_56 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c56
*+ bl_0_56 br_0_56 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c56
*+ bl_0_56 br_0_56 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c56
*+ bl_0_56 br_0_56 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c56
*+ bl_0_56 br_0_56 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c56
*+ bl_0_56 br_0_56 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c56
*+ bl_0_56 br_0_56 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c56
*+ bl_0_56 br_0_56 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c56
*+ bl_0_56 br_0_56 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c56
*+ bl_0_56 br_0_56 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c56
*+ bl_0_56 br_0_56 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c56
*+ bl_0_56 br_0_56 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c56
*+ bl_0_56 br_0_56 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c56
*+ bl_0_56 br_0_56 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c56
*+ bl_0_56 br_0_56 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c56
*+ bl_0_56 br_0_56 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c56
*+ bl_0_56 br_0_56 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c56
*+ bl_0_56 br_0_56 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c56
*+ bl_0_56 br_0_56 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c56
*+ bl_0_56 br_0_56 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c56
*+ bl_0_56 br_0_56 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c56
*+ bl_0_56 br_0_56 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c56
*+ bl_0_56 br_0_56 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c56
*+ bl_0_56 br_0_56 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c56
*+ bl_0_56 br_0_56 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c56
*+ bl_0_56 br_0_56 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c56
*+ bl_0_56 br_0_56 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c56
*+ bl_0_56 br_0_56 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c56
*+ bl_0_56 br_0_56 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c56
*+ bl_0_56 br_0_56 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c56
*+ bl_0_56 br_0_56 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c56
*+ bl_0_56 br_0_56 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c56
*+ bl_0_56 br_0_56 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c56
*+ bl_0_56 br_0_56 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c56
*+ bl_0_56 br_0_56 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c56
*+ bl_0_56 br_0_56 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c56
*+ bl_0_56 br_0_56 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c56
*+ bl_0_56 br_0_56 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c56
*+ bl_0_56 br_0_56 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c56
*+ bl_0_56 br_0_56 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c56
*+ bl_0_56 br_0_56 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c56
*+ bl_0_56 br_0_56 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c56
*+ bl_0_56 br_0_56 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c56
*+ bl_0_56 br_0_56 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c56
*+ bl_0_56 br_0_56 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c56
*+ bl_0_56 br_0_56 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c56
*+ bl_0_56 br_0_56 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c56
*+ bl_0_56 br_0_56 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c56
*+ bl_0_56 br_0_56 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c56
*+ bl_0_56 br_0_56 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c56
*+ bl_0_56 br_0_56 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c56
*+ bl_0_56 br_0_56 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c56
*+ bl_0_56 br_0_56 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c56
*+ bl_0_56 br_0_56 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c56
*+ bl_0_56 br_0_56 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c56
*+ bl_0_56 br_0_56 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c56
*+ bl_0_56 br_0_56 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c56
*+ bl_0_56 br_0_56 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c56
*+ bl_0_56 br_0_56 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c56
*+ bl_0_56 br_0_56 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c56
*+ bl_0_56 br_0_56 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c56
*+ bl_0_56 br_0_56 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c56
*+ bl_0_56 br_0_56 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c56
*+ bl_0_56 br_0_56 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c56
*+ bl_0_56 br_0_56 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c56
*+ bl_0_56 br_0_56 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c56
*+ bl_0_56 br_0_56 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c56
*+ bl_0_56 br_0_56 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c56
*+ bl_0_56 br_0_56 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c56
*+ bl_0_56 br_0_56 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c56
*+ bl_0_56 br_0_56 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c56
*+ bl_0_56 br_0_56 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c56
*+ bl_0_56 br_0_56 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c56
*+ bl_0_56 br_0_56 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c56
*+ bl_0_56 br_0_56 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c56
*+ bl_0_56 br_0_56 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c56
*+ bl_0_56 br_0_56 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c56
*+ bl_0_56 br_0_56 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c56
*+ bl_0_56 br_0_56 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c56
*+ bl_0_56 br_0_56 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c56
*+ bl_0_56 br_0_56 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c56
*+ bl_0_56 br_0_56 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c56
*+ bl_0_56 br_0_56 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c56
*+ bl_0_56 br_0_56 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c56
*+ bl_0_56 br_0_56 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c56
*+ bl_0_56 br_0_56 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c56
*+ bl_0_56 br_0_56 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c56
*+ bl_0_56 br_0_56 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c56
*+ bl_0_56 br_0_56 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c56
*+ bl_0_56 br_0_56 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c56
*+ bl_0_56 br_0_56 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c56
*+ bl_0_56 br_0_56 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c56
*+ bl_0_56 br_0_56 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c56
*+ bl_0_56 br_0_56 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c56
*+ bl_0_56 br_0_56 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c56
*+ bl_0_56 br_0_56 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c56
*+ bl_0_56 br_0_56 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c56
*+ bl_0_56 br_0_56 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c56
*+ bl_0_56 br_0_56 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c56
+ bl_0_56 br_0_56 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c57
+ bl_0_57 br_0_57 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c57
*+ bl_0_57 br_0_57 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c57
*+ bl_0_57 br_0_57 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c57
*+ bl_0_57 br_0_57 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c57
*+ bl_0_57 br_0_57 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c57
*+ bl_0_57 br_0_57 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c57
*+ bl_0_57 br_0_57 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c57
*+ bl_0_57 br_0_57 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c57
*+ bl_0_57 br_0_57 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c57
*+ bl_0_57 br_0_57 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c57
*+ bl_0_57 br_0_57 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c57
*+ bl_0_57 br_0_57 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c57
*+ bl_0_57 br_0_57 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c57
*+ bl_0_57 br_0_57 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c57
*+ bl_0_57 br_0_57 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c57
*+ bl_0_57 br_0_57 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c57
*+ bl_0_57 br_0_57 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c57
*+ bl_0_57 br_0_57 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c57
*+ bl_0_57 br_0_57 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c57
*+ bl_0_57 br_0_57 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c57
*+ bl_0_57 br_0_57 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c57
*+ bl_0_57 br_0_57 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c57
*+ bl_0_57 br_0_57 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c57
*+ bl_0_57 br_0_57 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c57
*+ bl_0_57 br_0_57 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c57
*+ bl_0_57 br_0_57 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c57
*+ bl_0_57 br_0_57 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c57
*+ bl_0_57 br_0_57 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c57
*+ bl_0_57 br_0_57 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c57
*+ bl_0_57 br_0_57 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c57
*+ bl_0_57 br_0_57 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c57
*+ bl_0_57 br_0_57 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c57
*+ bl_0_57 br_0_57 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c57
*+ bl_0_57 br_0_57 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c57
*+ bl_0_57 br_0_57 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c57
*+ bl_0_57 br_0_57 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c57
*+ bl_0_57 br_0_57 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c57
*+ bl_0_57 br_0_57 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c57
*+ bl_0_57 br_0_57 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c57
*+ bl_0_57 br_0_57 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c57
*+ bl_0_57 br_0_57 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c57
*+ bl_0_57 br_0_57 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c57
*+ bl_0_57 br_0_57 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c57
*+ bl_0_57 br_0_57 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c57
*+ bl_0_57 br_0_57 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c57
*+ bl_0_57 br_0_57 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c57
*+ bl_0_57 br_0_57 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c57
*+ bl_0_57 br_0_57 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c57
*+ bl_0_57 br_0_57 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c57
*+ bl_0_57 br_0_57 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c57
*+ bl_0_57 br_0_57 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c57
*+ bl_0_57 br_0_57 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c57
*+ bl_0_57 br_0_57 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c57
*+ bl_0_57 br_0_57 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c57
*+ bl_0_57 br_0_57 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c57
*+ bl_0_57 br_0_57 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c57
*+ bl_0_57 br_0_57 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c57
*+ bl_0_57 br_0_57 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c57
*+ bl_0_57 br_0_57 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c57
*+ bl_0_57 br_0_57 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c57
*+ bl_0_57 br_0_57 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c57
*+ bl_0_57 br_0_57 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c57
*+ bl_0_57 br_0_57 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c57
*+ bl_0_57 br_0_57 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c57
*+ bl_0_57 br_0_57 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c57
*+ bl_0_57 br_0_57 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c57
*+ bl_0_57 br_0_57 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c57
*+ bl_0_57 br_0_57 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c57
*+ bl_0_57 br_0_57 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c57
*+ bl_0_57 br_0_57 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c57
*+ bl_0_57 br_0_57 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c57
*+ bl_0_57 br_0_57 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c57
*+ bl_0_57 br_0_57 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c57
*+ bl_0_57 br_0_57 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c57
*+ bl_0_57 br_0_57 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c57
*+ bl_0_57 br_0_57 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c57
*+ bl_0_57 br_0_57 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c57
*+ bl_0_57 br_0_57 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c57
*+ bl_0_57 br_0_57 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c57
*+ bl_0_57 br_0_57 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c57
*+ bl_0_57 br_0_57 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c57
*+ bl_0_57 br_0_57 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c57
*+ bl_0_57 br_0_57 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c57
*+ bl_0_57 br_0_57 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c57
*+ bl_0_57 br_0_57 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c57
*+ bl_0_57 br_0_57 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c57
*+ bl_0_57 br_0_57 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c57
*+ bl_0_57 br_0_57 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c57
*+ bl_0_57 br_0_57 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c57
*+ bl_0_57 br_0_57 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c57
*+ bl_0_57 br_0_57 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c57
*+ bl_0_57 br_0_57 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c57
*+ bl_0_57 br_0_57 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c57
*+ bl_0_57 br_0_57 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c57
*+ bl_0_57 br_0_57 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c57
*+ bl_0_57 br_0_57 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c57
*+ bl_0_57 br_0_57 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c57
*+ bl_0_57 br_0_57 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c57
*+ bl_0_57 br_0_57 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c57
*+ bl_0_57 br_0_57 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c57
*+ bl_0_57 br_0_57 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c57
*+ bl_0_57 br_0_57 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c57
*+ bl_0_57 br_0_57 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c57
*+ bl_0_57 br_0_57 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c57
*+ bl_0_57 br_0_57 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c57
*+ bl_0_57 br_0_57 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c57
*+ bl_0_57 br_0_57 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c57
*+ bl_0_57 br_0_57 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c57
*+ bl_0_57 br_0_57 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c57
*+ bl_0_57 br_0_57 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c57
*+ bl_0_57 br_0_57 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c57
*+ bl_0_57 br_0_57 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c57
*+ bl_0_57 br_0_57 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c57
*+ bl_0_57 br_0_57 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c57
*+ bl_0_57 br_0_57 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c57
*+ bl_0_57 br_0_57 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c57
*+ bl_0_57 br_0_57 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c57
*+ bl_0_57 br_0_57 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c57
*+ bl_0_57 br_0_57 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c57
*+ bl_0_57 br_0_57 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c57
*+ bl_0_57 br_0_57 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c57
*+ bl_0_57 br_0_57 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c57
*+ bl_0_57 br_0_57 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c57
*+ bl_0_57 br_0_57 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c57
*+ bl_0_57 br_0_57 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c57
*+ bl_0_57 br_0_57 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c57
*+ bl_0_57 br_0_57 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c57
+ bl_0_57 br_0_57 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c58
+ bl_0_58 br_0_58 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c58
*+ bl_0_58 br_0_58 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c58
*+ bl_0_58 br_0_58 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c58
*+ bl_0_58 br_0_58 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c58
*+ bl_0_58 br_0_58 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c58
*+ bl_0_58 br_0_58 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c58
*+ bl_0_58 br_0_58 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c58
*+ bl_0_58 br_0_58 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c58
*+ bl_0_58 br_0_58 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c58
*+ bl_0_58 br_0_58 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c58
*+ bl_0_58 br_0_58 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c58
*+ bl_0_58 br_0_58 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c58
*+ bl_0_58 br_0_58 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c58
*+ bl_0_58 br_0_58 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c58
*+ bl_0_58 br_0_58 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c58
*+ bl_0_58 br_0_58 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c58
*+ bl_0_58 br_0_58 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c58
*+ bl_0_58 br_0_58 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c58
*+ bl_0_58 br_0_58 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c58
*+ bl_0_58 br_0_58 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c58
*+ bl_0_58 br_0_58 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c58
*+ bl_0_58 br_0_58 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c58
*+ bl_0_58 br_0_58 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c58
*+ bl_0_58 br_0_58 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c58
*+ bl_0_58 br_0_58 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c58
*+ bl_0_58 br_0_58 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c58
*+ bl_0_58 br_0_58 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c58
*+ bl_0_58 br_0_58 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c58
*+ bl_0_58 br_0_58 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c58
*+ bl_0_58 br_0_58 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c58
*+ bl_0_58 br_0_58 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c58
*+ bl_0_58 br_0_58 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c58
*+ bl_0_58 br_0_58 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c58
*+ bl_0_58 br_0_58 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c58
*+ bl_0_58 br_0_58 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c58
*+ bl_0_58 br_0_58 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c58
*+ bl_0_58 br_0_58 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c58
*+ bl_0_58 br_0_58 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c58
*+ bl_0_58 br_0_58 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c58
*+ bl_0_58 br_0_58 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c58
*+ bl_0_58 br_0_58 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c58
*+ bl_0_58 br_0_58 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c58
*+ bl_0_58 br_0_58 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c58
*+ bl_0_58 br_0_58 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c58
*+ bl_0_58 br_0_58 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c58
*+ bl_0_58 br_0_58 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c58
*+ bl_0_58 br_0_58 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c58
*+ bl_0_58 br_0_58 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c58
*+ bl_0_58 br_0_58 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c58
*+ bl_0_58 br_0_58 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c58
*+ bl_0_58 br_0_58 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c58
*+ bl_0_58 br_0_58 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c58
*+ bl_0_58 br_0_58 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c58
*+ bl_0_58 br_0_58 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c58
*+ bl_0_58 br_0_58 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c58
*+ bl_0_58 br_0_58 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c58
*+ bl_0_58 br_0_58 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c58
*+ bl_0_58 br_0_58 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c58
*+ bl_0_58 br_0_58 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c58
*+ bl_0_58 br_0_58 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c58
*+ bl_0_58 br_0_58 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c58
*+ bl_0_58 br_0_58 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c58
*+ bl_0_58 br_0_58 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c58
*+ bl_0_58 br_0_58 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c58
*+ bl_0_58 br_0_58 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c58
*+ bl_0_58 br_0_58 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c58
*+ bl_0_58 br_0_58 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c58
*+ bl_0_58 br_0_58 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c58
*+ bl_0_58 br_0_58 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c58
*+ bl_0_58 br_0_58 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c58
*+ bl_0_58 br_0_58 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c58
*+ bl_0_58 br_0_58 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c58
*+ bl_0_58 br_0_58 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c58
*+ bl_0_58 br_0_58 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c58
*+ bl_0_58 br_0_58 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c58
*+ bl_0_58 br_0_58 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c58
*+ bl_0_58 br_0_58 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c58
*+ bl_0_58 br_0_58 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c58
*+ bl_0_58 br_0_58 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c58
*+ bl_0_58 br_0_58 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c58
*+ bl_0_58 br_0_58 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c58
*+ bl_0_58 br_0_58 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c58
*+ bl_0_58 br_0_58 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c58
*+ bl_0_58 br_0_58 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c58
*+ bl_0_58 br_0_58 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c58
*+ bl_0_58 br_0_58 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c58
*+ bl_0_58 br_0_58 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c58
*+ bl_0_58 br_0_58 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c58
*+ bl_0_58 br_0_58 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c58
*+ bl_0_58 br_0_58 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c58
*+ bl_0_58 br_0_58 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c58
*+ bl_0_58 br_0_58 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c58
*+ bl_0_58 br_0_58 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c58
*+ bl_0_58 br_0_58 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c58
*+ bl_0_58 br_0_58 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c58
*+ bl_0_58 br_0_58 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c58
*+ bl_0_58 br_0_58 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c58
*+ bl_0_58 br_0_58 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c58
*+ bl_0_58 br_0_58 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c58
*+ bl_0_58 br_0_58 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c58
*+ bl_0_58 br_0_58 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c58
*+ bl_0_58 br_0_58 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c58
*+ bl_0_58 br_0_58 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c58
*+ bl_0_58 br_0_58 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c58
*+ bl_0_58 br_0_58 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c58
*+ bl_0_58 br_0_58 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c58
*+ bl_0_58 br_0_58 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c58
*+ bl_0_58 br_0_58 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c58
*+ bl_0_58 br_0_58 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c58
*+ bl_0_58 br_0_58 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c58
*+ bl_0_58 br_0_58 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c58
*+ bl_0_58 br_0_58 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c58
*+ bl_0_58 br_0_58 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c58
*+ bl_0_58 br_0_58 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c58
*+ bl_0_58 br_0_58 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c58
*+ bl_0_58 br_0_58 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c58
*+ bl_0_58 br_0_58 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c58
*+ bl_0_58 br_0_58 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c58
*+ bl_0_58 br_0_58 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c58
*+ bl_0_58 br_0_58 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c58
*+ bl_0_58 br_0_58 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c58
*+ bl_0_58 br_0_58 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c58
*+ bl_0_58 br_0_58 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c58
*+ bl_0_58 br_0_58 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c58
*+ bl_0_58 br_0_58 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c58
*+ bl_0_58 br_0_58 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c58
*+ bl_0_58 br_0_58 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c58
+ bl_0_58 br_0_58 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c59
+ bl_0_59 br_0_59 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c59
*+ bl_0_59 br_0_59 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c59
*+ bl_0_59 br_0_59 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c59
*+ bl_0_59 br_0_59 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c59
*+ bl_0_59 br_0_59 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c59
*+ bl_0_59 br_0_59 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c59
*+ bl_0_59 br_0_59 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c59
*+ bl_0_59 br_0_59 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c59
*+ bl_0_59 br_0_59 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c59
*+ bl_0_59 br_0_59 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c59
*+ bl_0_59 br_0_59 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c59
*+ bl_0_59 br_0_59 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c59
*+ bl_0_59 br_0_59 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c59
*+ bl_0_59 br_0_59 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c59
*+ bl_0_59 br_0_59 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c59
*+ bl_0_59 br_0_59 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c59
*+ bl_0_59 br_0_59 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c59
*+ bl_0_59 br_0_59 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c59
*+ bl_0_59 br_0_59 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c59
*+ bl_0_59 br_0_59 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c59
*+ bl_0_59 br_0_59 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c59
*+ bl_0_59 br_0_59 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c59
*+ bl_0_59 br_0_59 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c59
*+ bl_0_59 br_0_59 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c59
*+ bl_0_59 br_0_59 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c59
*+ bl_0_59 br_0_59 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c59
*+ bl_0_59 br_0_59 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c59
*+ bl_0_59 br_0_59 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c59
*+ bl_0_59 br_0_59 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c59
*+ bl_0_59 br_0_59 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c59
*+ bl_0_59 br_0_59 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c59
*+ bl_0_59 br_0_59 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c59
*+ bl_0_59 br_0_59 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c59
*+ bl_0_59 br_0_59 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c59
*+ bl_0_59 br_0_59 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c59
*+ bl_0_59 br_0_59 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c59
*+ bl_0_59 br_0_59 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c59
*+ bl_0_59 br_0_59 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c59
*+ bl_0_59 br_0_59 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c59
*+ bl_0_59 br_0_59 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c59
*+ bl_0_59 br_0_59 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c59
*+ bl_0_59 br_0_59 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c59
*+ bl_0_59 br_0_59 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c59
*+ bl_0_59 br_0_59 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c59
*+ bl_0_59 br_0_59 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c59
*+ bl_0_59 br_0_59 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c59
*+ bl_0_59 br_0_59 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c59
*+ bl_0_59 br_0_59 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c59
*+ bl_0_59 br_0_59 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c59
*+ bl_0_59 br_0_59 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c59
*+ bl_0_59 br_0_59 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c59
*+ bl_0_59 br_0_59 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c59
*+ bl_0_59 br_0_59 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c59
*+ bl_0_59 br_0_59 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c59
*+ bl_0_59 br_0_59 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c59
*+ bl_0_59 br_0_59 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c59
*+ bl_0_59 br_0_59 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c59
*+ bl_0_59 br_0_59 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c59
*+ bl_0_59 br_0_59 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c59
*+ bl_0_59 br_0_59 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c59
*+ bl_0_59 br_0_59 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c59
*+ bl_0_59 br_0_59 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c59
*+ bl_0_59 br_0_59 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c59
*+ bl_0_59 br_0_59 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c59
*+ bl_0_59 br_0_59 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c59
*+ bl_0_59 br_0_59 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c59
*+ bl_0_59 br_0_59 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c59
*+ bl_0_59 br_0_59 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c59
*+ bl_0_59 br_0_59 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c59
*+ bl_0_59 br_0_59 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c59
*+ bl_0_59 br_0_59 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c59
*+ bl_0_59 br_0_59 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c59
*+ bl_0_59 br_0_59 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c59
*+ bl_0_59 br_0_59 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c59
*+ bl_0_59 br_0_59 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c59
*+ bl_0_59 br_0_59 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c59
*+ bl_0_59 br_0_59 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c59
*+ bl_0_59 br_0_59 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c59
*+ bl_0_59 br_0_59 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c59
*+ bl_0_59 br_0_59 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c59
*+ bl_0_59 br_0_59 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c59
*+ bl_0_59 br_0_59 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c59
*+ bl_0_59 br_0_59 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c59
*+ bl_0_59 br_0_59 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c59
*+ bl_0_59 br_0_59 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c59
*+ bl_0_59 br_0_59 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c59
*+ bl_0_59 br_0_59 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c59
*+ bl_0_59 br_0_59 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c59
*+ bl_0_59 br_0_59 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c59
*+ bl_0_59 br_0_59 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c59
*+ bl_0_59 br_0_59 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c59
*+ bl_0_59 br_0_59 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c59
*+ bl_0_59 br_0_59 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c59
*+ bl_0_59 br_0_59 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c59
*+ bl_0_59 br_0_59 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c59
*+ bl_0_59 br_0_59 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c59
*+ bl_0_59 br_0_59 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c59
*+ bl_0_59 br_0_59 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c59
*+ bl_0_59 br_0_59 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c59
*+ bl_0_59 br_0_59 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c59
*+ bl_0_59 br_0_59 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c59
*+ bl_0_59 br_0_59 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c59
*+ bl_0_59 br_0_59 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c59
*+ bl_0_59 br_0_59 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c59
*+ bl_0_59 br_0_59 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c59
*+ bl_0_59 br_0_59 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c59
*+ bl_0_59 br_0_59 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c59
*+ bl_0_59 br_0_59 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c59
*+ bl_0_59 br_0_59 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c59
*+ bl_0_59 br_0_59 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c59
*+ bl_0_59 br_0_59 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c59
*+ bl_0_59 br_0_59 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c59
*+ bl_0_59 br_0_59 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c59
*+ bl_0_59 br_0_59 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c59
*+ bl_0_59 br_0_59 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c59
*+ bl_0_59 br_0_59 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c59
*+ bl_0_59 br_0_59 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c59
*+ bl_0_59 br_0_59 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c59
*+ bl_0_59 br_0_59 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c59
*+ bl_0_59 br_0_59 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c59
*+ bl_0_59 br_0_59 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c59
*+ bl_0_59 br_0_59 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c59
*+ bl_0_59 br_0_59 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c59
*+ bl_0_59 br_0_59 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c59
*+ bl_0_59 br_0_59 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c59
*+ bl_0_59 br_0_59 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c59
*+ bl_0_59 br_0_59 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c59
+ bl_0_59 br_0_59 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c60
+ bl_0_60 br_0_60 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c60
*+ bl_0_60 br_0_60 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c60
*+ bl_0_60 br_0_60 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c60
*+ bl_0_60 br_0_60 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c60
*+ bl_0_60 br_0_60 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c60
*+ bl_0_60 br_0_60 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c60
*+ bl_0_60 br_0_60 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c60
*+ bl_0_60 br_0_60 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c60
*+ bl_0_60 br_0_60 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c60
*+ bl_0_60 br_0_60 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c60
*+ bl_0_60 br_0_60 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c60
*+ bl_0_60 br_0_60 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c60
*+ bl_0_60 br_0_60 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c60
*+ bl_0_60 br_0_60 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c60
*+ bl_0_60 br_0_60 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c60
*+ bl_0_60 br_0_60 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c60
*+ bl_0_60 br_0_60 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c60
*+ bl_0_60 br_0_60 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c60
*+ bl_0_60 br_0_60 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c60
*+ bl_0_60 br_0_60 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c60
*+ bl_0_60 br_0_60 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c60
*+ bl_0_60 br_0_60 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c60
*+ bl_0_60 br_0_60 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c60
*+ bl_0_60 br_0_60 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c60
*+ bl_0_60 br_0_60 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c60
*+ bl_0_60 br_0_60 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c60
*+ bl_0_60 br_0_60 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c60
*+ bl_0_60 br_0_60 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c60
*+ bl_0_60 br_0_60 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c60
*+ bl_0_60 br_0_60 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c60
*+ bl_0_60 br_0_60 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c60
*+ bl_0_60 br_0_60 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c60
*+ bl_0_60 br_0_60 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c60
*+ bl_0_60 br_0_60 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c60
*+ bl_0_60 br_0_60 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c60
*+ bl_0_60 br_0_60 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c60
*+ bl_0_60 br_0_60 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c60
*+ bl_0_60 br_0_60 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c60
*+ bl_0_60 br_0_60 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c60
*+ bl_0_60 br_0_60 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c60
*+ bl_0_60 br_0_60 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c60
*+ bl_0_60 br_0_60 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c60
*+ bl_0_60 br_0_60 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c60
*+ bl_0_60 br_0_60 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c60
*+ bl_0_60 br_0_60 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c60
*+ bl_0_60 br_0_60 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c60
*+ bl_0_60 br_0_60 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c60
*+ bl_0_60 br_0_60 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c60
*+ bl_0_60 br_0_60 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c60
*+ bl_0_60 br_0_60 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c60
*+ bl_0_60 br_0_60 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c60
*+ bl_0_60 br_0_60 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c60
*+ bl_0_60 br_0_60 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c60
*+ bl_0_60 br_0_60 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c60
*+ bl_0_60 br_0_60 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c60
*+ bl_0_60 br_0_60 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c60
*+ bl_0_60 br_0_60 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c60
*+ bl_0_60 br_0_60 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c60
*+ bl_0_60 br_0_60 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c60
*+ bl_0_60 br_0_60 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c60
*+ bl_0_60 br_0_60 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c60
*+ bl_0_60 br_0_60 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c60
*+ bl_0_60 br_0_60 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c60
*+ bl_0_60 br_0_60 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c60
*+ bl_0_60 br_0_60 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c60
*+ bl_0_60 br_0_60 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c60
*+ bl_0_60 br_0_60 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c60
*+ bl_0_60 br_0_60 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c60
*+ bl_0_60 br_0_60 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c60
*+ bl_0_60 br_0_60 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c60
*+ bl_0_60 br_0_60 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c60
*+ bl_0_60 br_0_60 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c60
*+ bl_0_60 br_0_60 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c60
*+ bl_0_60 br_0_60 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c60
*+ bl_0_60 br_0_60 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c60
*+ bl_0_60 br_0_60 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c60
*+ bl_0_60 br_0_60 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c60
*+ bl_0_60 br_0_60 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c60
*+ bl_0_60 br_0_60 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c60
*+ bl_0_60 br_0_60 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c60
*+ bl_0_60 br_0_60 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c60
*+ bl_0_60 br_0_60 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c60
*+ bl_0_60 br_0_60 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c60
*+ bl_0_60 br_0_60 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c60
*+ bl_0_60 br_0_60 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c60
*+ bl_0_60 br_0_60 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c60
*+ bl_0_60 br_0_60 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c60
*+ bl_0_60 br_0_60 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c60
*+ bl_0_60 br_0_60 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c60
*+ bl_0_60 br_0_60 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c60
*+ bl_0_60 br_0_60 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c60
*+ bl_0_60 br_0_60 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c60
*+ bl_0_60 br_0_60 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c60
*+ bl_0_60 br_0_60 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c60
*+ bl_0_60 br_0_60 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c60
*+ bl_0_60 br_0_60 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c60
*+ bl_0_60 br_0_60 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c60
*+ bl_0_60 br_0_60 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c60
*+ bl_0_60 br_0_60 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c60
*+ bl_0_60 br_0_60 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c60
*+ bl_0_60 br_0_60 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c60
*+ bl_0_60 br_0_60 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c60
*+ bl_0_60 br_0_60 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c60
*+ bl_0_60 br_0_60 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c60
*+ bl_0_60 br_0_60 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c60
*+ bl_0_60 br_0_60 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c60
*+ bl_0_60 br_0_60 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c60
*+ bl_0_60 br_0_60 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c60
*+ bl_0_60 br_0_60 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c60
*+ bl_0_60 br_0_60 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c60
*+ bl_0_60 br_0_60 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c60
*+ bl_0_60 br_0_60 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c60
*+ bl_0_60 br_0_60 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c60
*+ bl_0_60 br_0_60 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c60
*+ bl_0_60 br_0_60 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c60
*+ bl_0_60 br_0_60 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c60
*+ bl_0_60 br_0_60 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c60
*+ bl_0_60 br_0_60 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c60
*+ bl_0_60 br_0_60 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c60
*+ bl_0_60 br_0_60 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c60
*+ bl_0_60 br_0_60 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c60
*+ bl_0_60 br_0_60 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c60
*+ bl_0_60 br_0_60 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c60
*+ bl_0_60 br_0_60 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c60
*+ bl_0_60 br_0_60 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c60
*+ bl_0_60 br_0_60 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c60
*+ bl_0_60 br_0_60 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c60
+ bl_0_60 br_0_60 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c61
+ bl_0_61 br_0_61 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c61
*+ bl_0_61 br_0_61 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c61
*+ bl_0_61 br_0_61 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c61
*+ bl_0_61 br_0_61 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c61
*+ bl_0_61 br_0_61 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c61
*+ bl_0_61 br_0_61 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c61
*+ bl_0_61 br_0_61 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c61
*+ bl_0_61 br_0_61 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c61
*+ bl_0_61 br_0_61 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c61
*+ bl_0_61 br_0_61 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c61
*+ bl_0_61 br_0_61 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c61
*+ bl_0_61 br_0_61 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c61
*+ bl_0_61 br_0_61 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c61
*+ bl_0_61 br_0_61 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c61
*+ bl_0_61 br_0_61 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c61
*+ bl_0_61 br_0_61 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c61
*+ bl_0_61 br_0_61 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c61
*+ bl_0_61 br_0_61 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c61
*+ bl_0_61 br_0_61 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c61
*+ bl_0_61 br_0_61 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c61
*+ bl_0_61 br_0_61 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c61
*+ bl_0_61 br_0_61 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c61
*+ bl_0_61 br_0_61 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c61
*+ bl_0_61 br_0_61 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c61
*+ bl_0_61 br_0_61 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c61
*+ bl_0_61 br_0_61 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c61
*+ bl_0_61 br_0_61 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c61
*+ bl_0_61 br_0_61 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c61
*+ bl_0_61 br_0_61 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c61
*+ bl_0_61 br_0_61 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c61
*+ bl_0_61 br_0_61 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c61
*+ bl_0_61 br_0_61 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c61
*+ bl_0_61 br_0_61 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c61
*+ bl_0_61 br_0_61 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c61
*+ bl_0_61 br_0_61 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c61
*+ bl_0_61 br_0_61 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c61
*+ bl_0_61 br_0_61 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c61
*+ bl_0_61 br_0_61 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c61
*+ bl_0_61 br_0_61 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c61
*+ bl_0_61 br_0_61 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c61
*+ bl_0_61 br_0_61 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c61
*+ bl_0_61 br_0_61 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c61
*+ bl_0_61 br_0_61 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c61
*+ bl_0_61 br_0_61 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c61
*+ bl_0_61 br_0_61 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c61
*+ bl_0_61 br_0_61 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c61
*+ bl_0_61 br_0_61 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c61
*+ bl_0_61 br_0_61 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c61
*+ bl_0_61 br_0_61 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c61
*+ bl_0_61 br_0_61 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c61
*+ bl_0_61 br_0_61 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c61
*+ bl_0_61 br_0_61 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c61
*+ bl_0_61 br_0_61 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c61
*+ bl_0_61 br_0_61 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c61
*+ bl_0_61 br_0_61 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c61
*+ bl_0_61 br_0_61 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c61
*+ bl_0_61 br_0_61 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c61
*+ bl_0_61 br_0_61 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c61
*+ bl_0_61 br_0_61 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c61
*+ bl_0_61 br_0_61 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c61
*+ bl_0_61 br_0_61 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c61
*+ bl_0_61 br_0_61 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c61
*+ bl_0_61 br_0_61 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c61
*+ bl_0_61 br_0_61 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c61
*+ bl_0_61 br_0_61 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c61
*+ bl_0_61 br_0_61 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c61
*+ bl_0_61 br_0_61 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c61
*+ bl_0_61 br_0_61 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c61
*+ bl_0_61 br_0_61 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c61
*+ bl_0_61 br_0_61 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c61
*+ bl_0_61 br_0_61 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c61
*+ bl_0_61 br_0_61 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c61
*+ bl_0_61 br_0_61 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c61
*+ bl_0_61 br_0_61 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c61
*+ bl_0_61 br_0_61 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c61
*+ bl_0_61 br_0_61 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c61
*+ bl_0_61 br_0_61 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c61
*+ bl_0_61 br_0_61 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c61
*+ bl_0_61 br_0_61 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c61
*+ bl_0_61 br_0_61 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c61
*+ bl_0_61 br_0_61 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c61
*+ bl_0_61 br_0_61 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c61
*+ bl_0_61 br_0_61 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c61
*+ bl_0_61 br_0_61 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c61
*+ bl_0_61 br_0_61 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c61
*+ bl_0_61 br_0_61 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c61
*+ bl_0_61 br_0_61 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c61
*+ bl_0_61 br_0_61 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c61
*+ bl_0_61 br_0_61 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c61
*+ bl_0_61 br_0_61 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c61
*+ bl_0_61 br_0_61 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c61
*+ bl_0_61 br_0_61 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c61
*+ bl_0_61 br_0_61 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c61
*+ bl_0_61 br_0_61 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c61
*+ bl_0_61 br_0_61 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c61
*+ bl_0_61 br_0_61 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c61
*+ bl_0_61 br_0_61 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c61
*+ bl_0_61 br_0_61 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c61
*+ bl_0_61 br_0_61 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c61
*+ bl_0_61 br_0_61 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c61
*+ bl_0_61 br_0_61 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c61
*+ bl_0_61 br_0_61 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c61
*+ bl_0_61 br_0_61 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c61
*+ bl_0_61 br_0_61 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c61
*+ bl_0_61 br_0_61 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c61
*+ bl_0_61 br_0_61 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c61
*+ bl_0_61 br_0_61 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c61
*+ bl_0_61 br_0_61 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c61
*+ bl_0_61 br_0_61 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c61
*+ bl_0_61 br_0_61 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c61
*+ bl_0_61 br_0_61 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c61
*+ bl_0_61 br_0_61 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c61
*+ bl_0_61 br_0_61 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c61
*+ bl_0_61 br_0_61 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c61
*+ bl_0_61 br_0_61 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c61
*+ bl_0_61 br_0_61 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c61
*+ bl_0_61 br_0_61 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c61
*+ bl_0_61 br_0_61 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c61
*+ bl_0_61 br_0_61 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c61
*+ bl_0_61 br_0_61 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c61
*+ bl_0_61 br_0_61 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c61
*+ bl_0_61 br_0_61 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c61
*+ bl_0_61 br_0_61 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c61
*+ bl_0_61 br_0_61 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c61
*+ bl_0_61 br_0_61 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c61
*+ bl_0_61 br_0_61 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c61
*+ bl_0_61 br_0_61 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c61
+ bl_0_61 br_0_61 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c62
+ bl_0_62 br_0_62 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c62
*+ bl_0_62 br_0_62 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c62
*+ bl_0_62 br_0_62 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c62
*+ bl_0_62 br_0_62 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c62
*+ bl_0_62 br_0_62 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c62
*+ bl_0_62 br_0_62 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c62
*+ bl_0_62 br_0_62 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c62
*+ bl_0_62 br_0_62 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c62
*+ bl_0_62 br_0_62 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c62
*+ bl_0_62 br_0_62 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c62
*+ bl_0_62 br_0_62 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c62
*+ bl_0_62 br_0_62 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c62
*+ bl_0_62 br_0_62 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c62
*+ bl_0_62 br_0_62 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c62
*+ bl_0_62 br_0_62 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c62
*+ bl_0_62 br_0_62 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c62
*+ bl_0_62 br_0_62 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c62
*+ bl_0_62 br_0_62 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c62
*+ bl_0_62 br_0_62 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c62
*+ bl_0_62 br_0_62 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c62
*+ bl_0_62 br_0_62 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c62
*+ bl_0_62 br_0_62 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c62
*+ bl_0_62 br_0_62 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c62
*+ bl_0_62 br_0_62 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c62
*+ bl_0_62 br_0_62 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c62
*+ bl_0_62 br_0_62 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c62
*+ bl_0_62 br_0_62 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c62
*+ bl_0_62 br_0_62 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c62
*+ bl_0_62 br_0_62 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c62
*+ bl_0_62 br_0_62 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c62
*+ bl_0_62 br_0_62 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c62
*+ bl_0_62 br_0_62 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c62
*+ bl_0_62 br_0_62 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c62
*+ bl_0_62 br_0_62 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c62
*+ bl_0_62 br_0_62 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c62
*+ bl_0_62 br_0_62 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c62
*+ bl_0_62 br_0_62 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c62
*+ bl_0_62 br_0_62 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c62
*+ bl_0_62 br_0_62 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c62
*+ bl_0_62 br_0_62 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c62
*+ bl_0_62 br_0_62 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c62
*+ bl_0_62 br_0_62 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c62
*+ bl_0_62 br_0_62 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c62
*+ bl_0_62 br_0_62 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c62
*+ bl_0_62 br_0_62 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c62
*+ bl_0_62 br_0_62 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c62
*+ bl_0_62 br_0_62 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c62
*+ bl_0_62 br_0_62 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c62
*+ bl_0_62 br_0_62 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c62
*+ bl_0_62 br_0_62 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c62
*+ bl_0_62 br_0_62 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c62
*+ bl_0_62 br_0_62 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c62
*+ bl_0_62 br_0_62 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c62
*+ bl_0_62 br_0_62 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c62
*+ bl_0_62 br_0_62 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c62
*+ bl_0_62 br_0_62 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c62
*+ bl_0_62 br_0_62 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c62
*+ bl_0_62 br_0_62 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c62
*+ bl_0_62 br_0_62 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c62
*+ bl_0_62 br_0_62 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c62
*+ bl_0_62 br_0_62 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c62
*+ bl_0_62 br_0_62 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c62
*+ bl_0_62 br_0_62 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c62
*+ bl_0_62 br_0_62 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c62
*+ bl_0_62 br_0_62 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c62
*+ bl_0_62 br_0_62 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c62
*+ bl_0_62 br_0_62 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c62
*+ bl_0_62 br_0_62 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c62
*+ bl_0_62 br_0_62 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c62
*+ bl_0_62 br_0_62 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c62
*+ bl_0_62 br_0_62 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c62
*+ bl_0_62 br_0_62 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c62
*+ bl_0_62 br_0_62 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c62
*+ bl_0_62 br_0_62 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c62
*+ bl_0_62 br_0_62 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c62
*+ bl_0_62 br_0_62 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c62
*+ bl_0_62 br_0_62 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c62
*+ bl_0_62 br_0_62 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c62
*+ bl_0_62 br_0_62 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c62
*+ bl_0_62 br_0_62 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c62
*+ bl_0_62 br_0_62 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c62
*+ bl_0_62 br_0_62 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c62
*+ bl_0_62 br_0_62 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c62
*+ bl_0_62 br_0_62 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c62
*+ bl_0_62 br_0_62 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c62
*+ bl_0_62 br_0_62 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c62
*+ bl_0_62 br_0_62 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c62
*+ bl_0_62 br_0_62 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c62
*+ bl_0_62 br_0_62 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c62
*+ bl_0_62 br_0_62 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c62
*+ bl_0_62 br_0_62 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c62
*+ bl_0_62 br_0_62 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c62
*+ bl_0_62 br_0_62 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c62
*+ bl_0_62 br_0_62 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c62
*+ bl_0_62 br_0_62 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c62
*+ bl_0_62 br_0_62 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c62
*+ bl_0_62 br_0_62 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c62
*+ bl_0_62 br_0_62 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c62
*+ bl_0_62 br_0_62 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c62
*+ bl_0_62 br_0_62 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c62
*+ bl_0_62 br_0_62 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c62
*+ bl_0_62 br_0_62 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c62
*+ bl_0_62 br_0_62 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c62
*+ bl_0_62 br_0_62 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c62
*+ bl_0_62 br_0_62 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c62
*+ bl_0_62 br_0_62 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c62
*+ bl_0_62 br_0_62 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c62
*+ bl_0_62 br_0_62 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c62
*+ bl_0_62 br_0_62 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c62
*+ bl_0_62 br_0_62 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c62
*+ bl_0_62 br_0_62 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c62
*+ bl_0_62 br_0_62 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c62
*+ bl_0_62 br_0_62 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c62
*+ bl_0_62 br_0_62 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c62
*+ bl_0_62 br_0_62 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c62
*+ bl_0_62 br_0_62 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c62
*+ bl_0_62 br_0_62 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c62
*+ bl_0_62 br_0_62 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c62
*+ bl_0_62 br_0_62 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c62
*+ bl_0_62 br_0_62 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c62
*+ bl_0_62 br_0_62 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c62
*+ bl_0_62 br_0_62 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c62
*+ bl_0_62 br_0_62 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c62
*+ bl_0_62 br_0_62 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c62
*+ bl_0_62 br_0_62 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c62
*+ bl_0_62 br_0_62 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c62
*+ bl_0_62 br_0_62 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c62
+ bl_0_62 br_0_62 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c63
+ bl_0_63 br_0_63 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c63
*+ bl_0_63 br_0_63 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c63
*+ bl_0_63 br_0_63 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c63
*+ bl_0_63 br_0_63 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c63
*+ bl_0_63 br_0_63 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c63
*+ bl_0_63 br_0_63 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c63
*+ bl_0_63 br_0_63 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c63
*+ bl_0_63 br_0_63 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c63
*+ bl_0_63 br_0_63 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c63
*+ bl_0_63 br_0_63 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c63
*+ bl_0_63 br_0_63 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c63
*+ bl_0_63 br_0_63 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c63
*+ bl_0_63 br_0_63 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c63
*+ bl_0_63 br_0_63 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c63
*+ bl_0_63 br_0_63 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c63
*+ bl_0_63 br_0_63 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c63
*+ bl_0_63 br_0_63 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c63
*+ bl_0_63 br_0_63 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c63
*+ bl_0_63 br_0_63 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c63
*+ bl_0_63 br_0_63 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c63
*+ bl_0_63 br_0_63 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c63
*+ bl_0_63 br_0_63 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c63
*+ bl_0_63 br_0_63 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c63
*+ bl_0_63 br_0_63 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c63
*+ bl_0_63 br_0_63 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c63
*+ bl_0_63 br_0_63 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c63
*+ bl_0_63 br_0_63 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c63
*+ bl_0_63 br_0_63 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c63
*+ bl_0_63 br_0_63 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c63
*+ bl_0_63 br_0_63 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c63
*+ bl_0_63 br_0_63 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c63
*+ bl_0_63 br_0_63 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c63
*+ bl_0_63 br_0_63 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c63
*+ bl_0_63 br_0_63 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c63
*+ bl_0_63 br_0_63 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c63
*+ bl_0_63 br_0_63 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c63
*+ bl_0_63 br_0_63 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c63
*+ bl_0_63 br_0_63 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c63
*+ bl_0_63 br_0_63 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c63
*+ bl_0_63 br_0_63 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c63
*+ bl_0_63 br_0_63 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c63
*+ bl_0_63 br_0_63 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c63
*+ bl_0_63 br_0_63 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c63
*+ bl_0_63 br_0_63 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c63
*+ bl_0_63 br_0_63 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c63
*+ bl_0_63 br_0_63 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c63
*+ bl_0_63 br_0_63 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c63
*+ bl_0_63 br_0_63 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c63
*+ bl_0_63 br_0_63 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c63
*+ bl_0_63 br_0_63 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c63
*+ bl_0_63 br_0_63 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c63
*+ bl_0_63 br_0_63 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c63
*+ bl_0_63 br_0_63 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c63
*+ bl_0_63 br_0_63 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c63
*+ bl_0_63 br_0_63 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c63
*+ bl_0_63 br_0_63 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c63
*+ bl_0_63 br_0_63 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c63
*+ bl_0_63 br_0_63 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c63
*+ bl_0_63 br_0_63 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c63
*+ bl_0_63 br_0_63 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c63
*+ bl_0_63 br_0_63 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c63
*+ bl_0_63 br_0_63 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c63
*+ bl_0_63 br_0_63 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c63
*+ bl_0_63 br_0_63 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c63
*+ bl_0_63 br_0_63 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c63
*+ bl_0_63 br_0_63 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c63
*+ bl_0_63 br_0_63 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c63
*+ bl_0_63 br_0_63 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c63
*+ bl_0_63 br_0_63 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c63
*+ bl_0_63 br_0_63 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c63
*+ bl_0_63 br_0_63 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c63
*+ bl_0_63 br_0_63 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c63
*+ bl_0_63 br_0_63 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c63
*+ bl_0_63 br_0_63 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c63
*+ bl_0_63 br_0_63 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c63
*+ bl_0_63 br_0_63 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c63
*+ bl_0_63 br_0_63 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c63
*+ bl_0_63 br_0_63 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c63
*+ bl_0_63 br_0_63 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c63
*+ bl_0_63 br_0_63 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c63
*+ bl_0_63 br_0_63 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c63
*+ bl_0_63 br_0_63 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c63
*+ bl_0_63 br_0_63 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c63
*+ bl_0_63 br_0_63 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c63
*+ bl_0_63 br_0_63 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c63
*+ bl_0_63 br_0_63 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c63
*+ bl_0_63 br_0_63 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c63
*+ bl_0_63 br_0_63 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c63
*+ bl_0_63 br_0_63 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c63
*+ bl_0_63 br_0_63 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c63
*+ bl_0_63 br_0_63 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c63
*+ bl_0_63 br_0_63 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c63
*+ bl_0_63 br_0_63 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c63
*+ bl_0_63 br_0_63 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c63
*+ bl_0_63 br_0_63 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c63
*+ bl_0_63 br_0_63 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c63
*+ bl_0_63 br_0_63 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c63
*+ bl_0_63 br_0_63 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c63
*+ bl_0_63 br_0_63 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c63
*+ bl_0_63 br_0_63 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c63
*+ bl_0_63 br_0_63 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c63
*+ bl_0_63 br_0_63 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c63
*+ bl_0_63 br_0_63 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c63
*+ bl_0_63 br_0_63 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c63
*+ bl_0_63 br_0_63 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c63
*+ bl_0_63 br_0_63 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c63
*+ bl_0_63 br_0_63 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c63
*+ bl_0_63 br_0_63 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c63
*+ bl_0_63 br_0_63 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c63
*+ bl_0_63 br_0_63 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c63
*+ bl_0_63 br_0_63 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c63
*+ bl_0_63 br_0_63 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c63
*+ bl_0_63 br_0_63 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c63
*+ bl_0_63 br_0_63 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c63
*+ bl_0_63 br_0_63 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c63
*+ bl_0_63 br_0_63 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c63
*+ bl_0_63 br_0_63 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c63
*+ bl_0_63 br_0_63 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c63
*+ bl_0_63 br_0_63 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c63
*+ bl_0_63 br_0_63 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c63
*+ bl_0_63 br_0_63 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c63
*+ bl_0_63 br_0_63 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c63
*+ bl_0_63 br_0_63 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c63
*+ bl_0_63 br_0_63 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c63
*+ bl_0_63 br_0_63 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c63
*+ bl_0_63 br_0_63 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c63
*+ bl_0_63 br_0_63 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c63
+ bl_0_63 br_0_63 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c64
+ bl_0_64 br_0_64 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c64
*+ bl_0_64 br_0_64 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c64
*+ bl_0_64 br_0_64 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c64
*+ bl_0_64 br_0_64 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c64
*+ bl_0_64 br_0_64 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c64
*+ bl_0_64 br_0_64 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c64
*+ bl_0_64 br_0_64 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c64
*+ bl_0_64 br_0_64 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c64
*+ bl_0_64 br_0_64 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c64
*+ bl_0_64 br_0_64 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c64
*+ bl_0_64 br_0_64 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c64
*+ bl_0_64 br_0_64 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c64
*+ bl_0_64 br_0_64 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c64
*+ bl_0_64 br_0_64 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c64
*+ bl_0_64 br_0_64 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c64
*+ bl_0_64 br_0_64 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c64
*+ bl_0_64 br_0_64 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c64
*+ bl_0_64 br_0_64 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c64
*+ bl_0_64 br_0_64 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c64
*+ bl_0_64 br_0_64 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c64
*+ bl_0_64 br_0_64 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c64
*+ bl_0_64 br_0_64 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c64
*+ bl_0_64 br_0_64 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c64
*+ bl_0_64 br_0_64 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c64
*+ bl_0_64 br_0_64 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c64
*+ bl_0_64 br_0_64 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c64
*+ bl_0_64 br_0_64 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c64
*+ bl_0_64 br_0_64 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c64
*+ bl_0_64 br_0_64 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c64
*+ bl_0_64 br_0_64 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c64
*+ bl_0_64 br_0_64 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c64
*+ bl_0_64 br_0_64 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c64
*+ bl_0_64 br_0_64 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c64
*+ bl_0_64 br_0_64 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c64
*+ bl_0_64 br_0_64 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c64
*+ bl_0_64 br_0_64 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c64
*+ bl_0_64 br_0_64 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c64
*+ bl_0_64 br_0_64 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c64
*+ bl_0_64 br_0_64 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c64
*+ bl_0_64 br_0_64 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c64
*+ bl_0_64 br_0_64 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c64
*+ bl_0_64 br_0_64 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c64
*+ bl_0_64 br_0_64 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c64
*+ bl_0_64 br_0_64 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c64
*+ bl_0_64 br_0_64 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c64
*+ bl_0_64 br_0_64 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c64
*+ bl_0_64 br_0_64 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c64
*+ bl_0_64 br_0_64 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c64
*+ bl_0_64 br_0_64 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c64
*+ bl_0_64 br_0_64 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c64
*+ bl_0_64 br_0_64 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c64
*+ bl_0_64 br_0_64 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c64
*+ bl_0_64 br_0_64 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c64
*+ bl_0_64 br_0_64 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c64
*+ bl_0_64 br_0_64 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c64
*+ bl_0_64 br_0_64 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c64
*+ bl_0_64 br_0_64 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c64
*+ bl_0_64 br_0_64 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c64
*+ bl_0_64 br_0_64 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c64
*+ bl_0_64 br_0_64 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c64
*+ bl_0_64 br_0_64 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c64
*+ bl_0_64 br_0_64 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c64
*+ bl_0_64 br_0_64 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c64
*+ bl_0_64 br_0_64 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c64
*+ bl_0_64 br_0_64 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c64
*+ bl_0_64 br_0_64 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c64
*+ bl_0_64 br_0_64 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c64
*+ bl_0_64 br_0_64 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c64
*+ bl_0_64 br_0_64 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c64
*+ bl_0_64 br_0_64 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c64
*+ bl_0_64 br_0_64 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c64
*+ bl_0_64 br_0_64 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c64
*+ bl_0_64 br_0_64 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c64
*+ bl_0_64 br_0_64 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c64
*+ bl_0_64 br_0_64 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c64
*+ bl_0_64 br_0_64 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c64
*+ bl_0_64 br_0_64 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c64
*+ bl_0_64 br_0_64 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c64
*+ bl_0_64 br_0_64 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c64
*+ bl_0_64 br_0_64 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c64
*+ bl_0_64 br_0_64 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c64
*+ bl_0_64 br_0_64 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c64
*+ bl_0_64 br_0_64 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c64
*+ bl_0_64 br_0_64 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c64
*+ bl_0_64 br_0_64 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c64
*+ bl_0_64 br_0_64 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c64
*+ bl_0_64 br_0_64 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c64
*+ bl_0_64 br_0_64 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c64
*+ bl_0_64 br_0_64 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c64
*+ bl_0_64 br_0_64 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c64
*+ bl_0_64 br_0_64 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c64
*+ bl_0_64 br_0_64 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c64
*+ bl_0_64 br_0_64 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c64
*+ bl_0_64 br_0_64 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c64
*+ bl_0_64 br_0_64 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c64
*+ bl_0_64 br_0_64 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c64
*+ bl_0_64 br_0_64 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c64
*+ bl_0_64 br_0_64 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c64
*+ bl_0_64 br_0_64 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c64
*+ bl_0_64 br_0_64 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c64
*+ bl_0_64 br_0_64 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c64
*+ bl_0_64 br_0_64 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c64
*+ bl_0_64 br_0_64 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c64
*+ bl_0_64 br_0_64 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c64
*+ bl_0_64 br_0_64 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c64
*+ bl_0_64 br_0_64 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c64
*+ bl_0_64 br_0_64 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c64
*+ bl_0_64 br_0_64 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c64
*+ bl_0_64 br_0_64 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c64
*+ bl_0_64 br_0_64 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c64
*+ bl_0_64 br_0_64 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c64
*+ bl_0_64 br_0_64 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c64
*+ bl_0_64 br_0_64 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c64
*+ bl_0_64 br_0_64 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c64
*+ bl_0_64 br_0_64 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c64
*+ bl_0_64 br_0_64 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c64
*+ bl_0_64 br_0_64 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c64
*+ bl_0_64 br_0_64 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c64
*+ bl_0_64 br_0_64 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c64
*+ bl_0_64 br_0_64 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c64
*+ bl_0_64 br_0_64 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c64
*+ bl_0_64 br_0_64 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c64
*+ bl_0_64 br_0_64 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c64
*+ bl_0_64 br_0_64 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c64
*+ bl_0_64 br_0_64 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c64
*+ bl_0_64 br_0_64 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c64
*+ bl_0_64 br_0_64 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c64
+ bl_0_64 br_0_64 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c65
+ bl_0_65 br_0_65 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c65
*+ bl_0_65 br_0_65 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c65
*+ bl_0_65 br_0_65 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c65
*+ bl_0_65 br_0_65 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c65
*+ bl_0_65 br_0_65 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c65
*+ bl_0_65 br_0_65 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c65
*+ bl_0_65 br_0_65 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c65
*+ bl_0_65 br_0_65 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c65
*+ bl_0_65 br_0_65 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c65
*+ bl_0_65 br_0_65 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c65
*+ bl_0_65 br_0_65 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c65
*+ bl_0_65 br_0_65 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c65
*+ bl_0_65 br_0_65 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c65
*+ bl_0_65 br_0_65 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c65
*+ bl_0_65 br_0_65 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c65
*+ bl_0_65 br_0_65 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c65
*+ bl_0_65 br_0_65 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c65
*+ bl_0_65 br_0_65 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c65
*+ bl_0_65 br_0_65 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c65
*+ bl_0_65 br_0_65 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c65
*+ bl_0_65 br_0_65 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c65
*+ bl_0_65 br_0_65 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c65
*+ bl_0_65 br_0_65 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c65
*+ bl_0_65 br_0_65 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c65
*+ bl_0_65 br_0_65 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c65
*+ bl_0_65 br_0_65 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c65
*+ bl_0_65 br_0_65 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c65
*+ bl_0_65 br_0_65 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c65
*+ bl_0_65 br_0_65 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c65
*+ bl_0_65 br_0_65 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c65
*+ bl_0_65 br_0_65 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c65
*+ bl_0_65 br_0_65 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c65
*+ bl_0_65 br_0_65 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c65
*+ bl_0_65 br_0_65 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c65
*+ bl_0_65 br_0_65 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c65
*+ bl_0_65 br_0_65 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c65
*+ bl_0_65 br_0_65 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c65
*+ bl_0_65 br_0_65 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c65
*+ bl_0_65 br_0_65 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c65
*+ bl_0_65 br_0_65 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c65
*+ bl_0_65 br_0_65 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c65
*+ bl_0_65 br_0_65 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c65
*+ bl_0_65 br_0_65 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c65
*+ bl_0_65 br_0_65 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c65
*+ bl_0_65 br_0_65 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c65
*+ bl_0_65 br_0_65 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c65
*+ bl_0_65 br_0_65 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c65
*+ bl_0_65 br_0_65 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c65
*+ bl_0_65 br_0_65 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c65
*+ bl_0_65 br_0_65 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c65
*+ bl_0_65 br_0_65 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c65
*+ bl_0_65 br_0_65 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c65
*+ bl_0_65 br_0_65 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c65
*+ bl_0_65 br_0_65 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c65
*+ bl_0_65 br_0_65 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c65
*+ bl_0_65 br_0_65 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c65
*+ bl_0_65 br_0_65 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c65
*+ bl_0_65 br_0_65 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c65
*+ bl_0_65 br_0_65 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c65
*+ bl_0_65 br_0_65 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c65
*+ bl_0_65 br_0_65 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c65
*+ bl_0_65 br_0_65 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c65
*+ bl_0_65 br_0_65 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c65
*+ bl_0_65 br_0_65 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c65
*+ bl_0_65 br_0_65 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c65
*+ bl_0_65 br_0_65 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c65
*+ bl_0_65 br_0_65 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c65
*+ bl_0_65 br_0_65 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c65
*+ bl_0_65 br_0_65 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c65
*+ bl_0_65 br_0_65 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c65
*+ bl_0_65 br_0_65 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c65
*+ bl_0_65 br_0_65 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c65
*+ bl_0_65 br_0_65 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c65
*+ bl_0_65 br_0_65 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c65
*+ bl_0_65 br_0_65 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c65
*+ bl_0_65 br_0_65 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c65
*+ bl_0_65 br_0_65 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c65
*+ bl_0_65 br_0_65 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c65
*+ bl_0_65 br_0_65 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c65
*+ bl_0_65 br_0_65 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c65
*+ bl_0_65 br_0_65 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c65
*+ bl_0_65 br_0_65 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c65
*+ bl_0_65 br_0_65 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c65
*+ bl_0_65 br_0_65 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c65
*+ bl_0_65 br_0_65 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c65
*+ bl_0_65 br_0_65 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c65
*+ bl_0_65 br_0_65 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c65
*+ bl_0_65 br_0_65 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c65
*+ bl_0_65 br_0_65 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c65
*+ bl_0_65 br_0_65 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c65
*+ bl_0_65 br_0_65 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c65
*+ bl_0_65 br_0_65 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c65
*+ bl_0_65 br_0_65 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c65
*+ bl_0_65 br_0_65 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c65
*+ bl_0_65 br_0_65 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c65
*+ bl_0_65 br_0_65 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c65
*+ bl_0_65 br_0_65 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c65
*+ bl_0_65 br_0_65 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c65
*+ bl_0_65 br_0_65 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c65
*+ bl_0_65 br_0_65 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c65
*+ bl_0_65 br_0_65 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c65
*+ bl_0_65 br_0_65 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c65
*+ bl_0_65 br_0_65 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c65
*+ bl_0_65 br_0_65 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c65
*+ bl_0_65 br_0_65 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c65
*+ bl_0_65 br_0_65 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c65
*+ bl_0_65 br_0_65 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c65
*+ bl_0_65 br_0_65 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c65
*+ bl_0_65 br_0_65 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c65
*+ bl_0_65 br_0_65 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c65
*+ bl_0_65 br_0_65 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c65
*+ bl_0_65 br_0_65 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c65
*+ bl_0_65 br_0_65 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c65
*+ bl_0_65 br_0_65 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c65
*+ bl_0_65 br_0_65 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c65
*+ bl_0_65 br_0_65 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c65
*+ bl_0_65 br_0_65 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c65
*+ bl_0_65 br_0_65 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c65
*+ bl_0_65 br_0_65 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c65
*+ bl_0_65 br_0_65 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c65
*+ bl_0_65 br_0_65 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c65
*+ bl_0_65 br_0_65 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c65
*+ bl_0_65 br_0_65 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c65
*+ bl_0_65 br_0_65 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c65
*+ bl_0_65 br_0_65 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c65
*+ bl_0_65 br_0_65 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c65
*+ bl_0_65 br_0_65 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c65
+ bl_0_65 br_0_65 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c66
+ bl_0_66 br_0_66 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c66
*+ bl_0_66 br_0_66 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c66
*+ bl_0_66 br_0_66 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c66
*+ bl_0_66 br_0_66 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c66
*+ bl_0_66 br_0_66 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c66
*+ bl_0_66 br_0_66 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c66
*+ bl_0_66 br_0_66 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c66
*+ bl_0_66 br_0_66 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c66
*+ bl_0_66 br_0_66 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c66
*+ bl_0_66 br_0_66 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c66
*+ bl_0_66 br_0_66 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c66
*+ bl_0_66 br_0_66 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c66
*+ bl_0_66 br_0_66 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c66
*+ bl_0_66 br_0_66 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c66
*+ bl_0_66 br_0_66 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c66
*+ bl_0_66 br_0_66 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c66
*+ bl_0_66 br_0_66 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c66
*+ bl_0_66 br_0_66 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c66
*+ bl_0_66 br_0_66 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c66
*+ bl_0_66 br_0_66 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c66
*+ bl_0_66 br_0_66 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c66
*+ bl_0_66 br_0_66 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c66
*+ bl_0_66 br_0_66 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c66
*+ bl_0_66 br_0_66 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c66
*+ bl_0_66 br_0_66 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c66
*+ bl_0_66 br_0_66 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c66
*+ bl_0_66 br_0_66 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c66
*+ bl_0_66 br_0_66 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c66
*+ bl_0_66 br_0_66 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c66
*+ bl_0_66 br_0_66 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c66
*+ bl_0_66 br_0_66 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c66
*+ bl_0_66 br_0_66 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c66
*+ bl_0_66 br_0_66 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c66
*+ bl_0_66 br_0_66 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c66
*+ bl_0_66 br_0_66 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c66
*+ bl_0_66 br_0_66 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c66
*+ bl_0_66 br_0_66 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c66
*+ bl_0_66 br_0_66 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c66
*+ bl_0_66 br_0_66 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c66
*+ bl_0_66 br_0_66 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c66
*+ bl_0_66 br_0_66 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c66
*+ bl_0_66 br_0_66 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c66
*+ bl_0_66 br_0_66 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c66
*+ bl_0_66 br_0_66 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c66
*+ bl_0_66 br_0_66 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c66
*+ bl_0_66 br_0_66 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c66
*+ bl_0_66 br_0_66 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c66
*+ bl_0_66 br_0_66 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c66
*+ bl_0_66 br_0_66 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c66
*+ bl_0_66 br_0_66 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c66
*+ bl_0_66 br_0_66 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c66
*+ bl_0_66 br_0_66 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c66
*+ bl_0_66 br_0_66 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c66
*+ bl_0_66 br_0_66 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c66
*+ bl_0_66 br_0_66 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c66
*+ bl_0_66 br_0_66 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c66
*+ bl_0_66 br_0_66 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c66
*+ bl_0_66 br_0_66 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c66
*+ bl_0_66 br_0_66 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c66
*+ bl_0_66 br_0_66 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c66
*+ bl_0_66 br_0_66 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c66
*+ bl_0_66 br_0_66 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c66
*+ bl_0_66 br_0_66 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c66
*+ bl_0_66 br_0_66 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c66
*+ bl_0_66 br_0_66 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c66
*+ bl_0_66 br_0_66 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c66
*+ bl_0_66 br_0_66 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c66
*+ bl_0_66 br_0_66 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c66
*+ bl_0_66 br_0_66 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c66
*+ bl_0_66 br_0_66 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c66
*+ bl_0_66 br_0_66 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c66
*+ bl_0_66 br_0_66 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c66
*+ bl_0_66 br_0_66 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c66
*+ bl_0_66 br_0_66 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c66
*+ bl_0_66 br_0_66 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c66
*+ bl_0_66 br_0_66 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c66
*+ bl_0_66 br_0_66 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c66
*+ bl_0_66 br_0_66 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c66
*+ bl_0_66 br_0_66 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c66
*+ bl_0_66 br_0_66 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c66
*+ bl_0_66 br_0_66 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c66
*+ bl_0_66 br_0_66 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c66
*+ bl_0_66 br_0_66 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c66
*+ bl_0_66 br_0_66 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c66
*+ bl_0_66 br_0_66 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c66
*+ bl_0_66 br_0_66 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c66
*+ bl_0_66 br_0_66 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c66
*+ bl_0_66 br_0_66 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c66
*+ bl_0_66 br_0_66 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c66
*+ bl_0_66 br_0_66 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c66
*+ bl_0_66 br_0_66 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c66
*+ bl_0_66 br_0_66 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c66
*+ bl_0_66 br_0_66 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c66
*+ bl_0_66 br_0_66 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c66
*+ bl_0_66 br_0_66 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c66
*+ bl_0_66 br_0_66 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c66
*+ bl_0_66 br_0_66 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c66
*+ bl_0_66 br_0_66 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c66
*+ bl_0_66 br_0_66 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c66
*+ bl_0_66 br_0_66 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c66
*+ bl_0_66 br_0_66 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c66
*+ bl_0_66 br_0_66 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c66
*+ bl_0_66 br_0_66 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c66
*+ bl_0_66 br_0_66 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c66
*+ bl_0_66 br_0_66 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c66
*+ bl_0_66 br_0_66 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c66
*+ bl_0_66 br_0_66 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c66
*+ bl_0_66 br_0_66 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c66
*+ bl_0_66 br_0_66 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c66
*+ bl_0_66 br_0_66 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c66
*+ bl_0_66 br_0_66 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c66
*+ bl_0_66 br_0_66 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c66
*+ bl_0_66 br_0_66 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c66
*+ bl_0_66 br_0_66 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c66
*+ bl_0_66 br_0_66 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c66
*+ bl_0_66 br_0_66 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c66
*+ bl_0_66 br_0_66 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c66
*+ bl_0_66 br_0_66 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c66
*+ bl_0_66 br_0_66 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c66
*+ bl_0_66 br_0_66 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c66
*+ bl_0_66 br_0_66 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c66
*+ bl_0_66 br_0_66 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c66
*+ bl_0_66 br_0_66 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c66
*+ bl_0_66 br_0_66 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c66
*+ bl_0_66 br_0_66 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c66
*+ bl_0_66 br_0_66 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c66
*+ bl_0_66 br_0_66 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c66
+ bl_0_66 br_0_66 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c67
+ bl_0_67 br_0_67 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c67
*+ bl_0_67 br_0_67 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c67
*+ bl_0_67 br_0_67 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c67
*+ bl_0_67 br_0_67 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c67
*+ bl_0_67 br_0_67 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c67
*+ bl_0_67 br_0_67 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c67
*+ bl_0_67 br_0_67 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c67
*+ bl_0_67 br_0_67 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c67
*+ bl_0_67 br_0_67 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c67
*+ bl_0_67 br_0_67 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c67
*+ bl_0_67 br_0_67 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c67
*+ bl_0_67 br_0_67 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c67
*+ bl_0_67 br_0_67 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c67
*+ bl_0_67 br_0_67 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c67
*+ bl_0_67 br_0_67 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c67
*+ bl_0_67 br_0_67 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c67
*+ bl_0_67 br_0_67 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c67
*+ bl_0_67 br_0_67 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c67
*+ bl_0_67 br_0_67 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c67
*+ bl_0_67 br_0_67 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c67
*+ bl_0_67 br_0_67 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c67
*+ bl_0_67 br_0_67 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c67
*+ bl_0_67 br_0_67 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c67
*+ bl_0_67 br_0_67 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c67
*+ bl_0_67 br_0_67 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c67
*+ bl_0_67 br_0_67 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c67
*+ bl_0_67 br_0_67 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c67
*+ bl_0_67 br_0_67 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c67
*+ bl_0_67 br_0_67 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c67
*+ bl_0_67 br_0_67 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c67
*+ bl_0_67 br_0_67 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c67
*+ bl_0_67 br_0_67 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c67
*+ bl_0_67 br_0_67 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c67
*+ bl_0_67 br_0_67 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c67
*+ bl_0_67 br_0_67 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c67
*+ bl_0_67 br_0_67 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c67
*+ bl_0_67 br_0_67 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c67
*+ bl_0_67 br_0_67 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c67
*+ bl_0_67 br_0_67 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c67
*+ bl_0_67 br_0_67 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c67
*+ bl_0_67 br_0_67 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c67
*+ bl_0_67 br_0_67 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c67
*+ bl_0_67 br_0_67 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c67
*+ bl_0_67 br_0_67 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c67
*+ bl_0_67 br_0_67 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c67
*+ bl_0_67 br_0_67 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c67
*+ bl_0_67 br_0_67 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c67
*+ bl_0_67 br_0_67 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c67
*+ bl_0_67 br_0_67 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c67
*+ bl_0_67 br_0_67 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c67
*+ bl_0_67 br_0_67 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c67
*+ bl_0_67 br_0_67 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c67
*+ bl_0_67 br_0_67 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c67
*+ bl_0_67 br_0_67 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c67
*+ bl_0_67 br_0_67 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c67
*+ bl_0_67 br_0_67 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c67
*+ bl_0_67 br_0_67 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c67
*+ bl_0_67 br_0_67 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c67
*+ bl_0_67 br_0_67 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c67
*+ bl_0_67 br_0_67 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c67
*+ bl_0_67 br_0_67 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c67
*+ bl_0_67 br_0_67 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c67
*+ bl_0_67 br_0_67 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c67
*+ bl_0_67 br_0_67 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c67
*+ bl_0_67 br_0_67 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c67
*+ bl_0_67 br_0_67 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c67
*+ bl_0_67 br_0_67 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c67
*+ bl_0_67 br_0_67 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c67
*+ bl_0_67 br_0_67 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c67
*+ bl_0_67 br_0_67 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c67
*+ bl_0_67 br_0_67 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c67
*+ bl_0_67 br_0_67 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c67
*+ bl_0_67 br_0_67 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c67
*+ bl_0_67 br_0_67 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c67
*+ bl_0_67 br_0_67 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c67
*+ bl_0_67 br_0_67 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c67
*+ bl_0_67 br_0_67 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c67
*+ bl_0_67 br_0_67 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c67
*+ bl_0_67 br_0_67 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c67
*+ bl_0_67 br_0_67 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c67
*+ bl_0_67 br_0_67 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c67
*+ bl_0_67 br_0_67 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c67
*+ bl_0_67 br_0_67 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c67
*+ bl_0_67 br_0_67 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c67
*+ bl_0_67 br_0_67 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c67
*+ bl_0_67 br_0_67 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c67
*+ bl_0_67 br_0_67 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c67
*+ bl_0_67 br_0_67 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c67
*+ bl_0_67 br_0_67 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c67
*+ bl_0_67 br_0_67 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c67
*+ bl_0_67 br_0_67 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c67
*+ bl_0_67 br_0_67 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c67
*+ bl_0_67 br_0_67 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c67
*+ bl_0_67 br_0_67 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c67
*+ bl_0_67 br_0_67 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c67
*+ bl_0_67 br_0_67 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c67
*+ bl_0_67 br_0_67 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c67
*+ bl_0_67 br_0_67 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c67
*+ bl_0_67 br_0_67 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c67
*+ bl_0_67 br_0_67 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c67
*+ bl_0_67 br_0_67 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c67
*+ bl_0_67 br_0_67 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c67
*+ bl_0_67 br_0_67 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c67
*+ bl_0_67 br_0_67 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c67
*+ bl_0_67 br_0_67 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c67
*+ bl_0_67 br_0_67 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c67
*+ bl_0_67 br_0_67 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c67
*+ bl_0_67 br_0_67 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c67
*+ bl_0_67 br_0_67 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c67
*+ bl_0_67 br_0_67 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c67
*+ bl_0_67 br_0_67 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c67
*+ bl_0_67 br_0_67 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c67
*+ bl_0_67 br_0_67 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c67
*+ bl_0_67 br_0_67 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c67
*+ bl_0_67 br_0_67 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c67
*+ bl_0_67 br_0_67 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c67
*+ bl_0_67 br_0_67 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c67
*+ bl_0_67 br_0_67 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c67
*+ bl_0_67 br_0_67 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c67
*+ bl_0_67 br_0_67 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c67
*+ bl_0_67 br_0_67 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c67
*+ bl_0_67 br_0_67 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c67
*+ bl_0_67 br_0_67 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c67
*+ bl_0_67 br_0_67 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c67
*+ bl_0_67 br_0_67 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c67
*+ bl_0_67 br_0_67 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c67
*+ bl_0_67 br_0_67 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c67
+ bl_0_67 br_0_67 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c68
+ bl_0_68 br_0_68 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c68
*+ bl_0_68 br_0_68 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c68
*+ bl_0_68 br_0_68 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c68
*+ bl_0_68 br_0_68 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c68
*+ bl_0_68 br_0_68 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c68
*+ bl_0_68 br_0_68 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c68
*+ bl_0_68 br_0_68 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c68
*+ bl_0_68 br_0_68 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c68
*+ bl_0_68 br_0_68 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c68
*+ bl_0_68 br_0_68 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c68
*+ bl_0_68 br_0_68 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c68
*+ bl_0_68 br_0_68 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c68
*+ bl_0_68 br_0_68 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c68
*+ bl_0_68 br_0_68 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c68
*+ bl_0_68 br_0_68 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c68
*+ bl_0_68 br_0_68 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c68
*+ bl_0_68 br_0_68 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c68
*+ bl_0_68 br_0_68 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c68
*+ bl_0_68 br_0_68 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c68
*+ bl_0_68 br_0_68 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c68
*+ bl_0_68 br_0_68 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c68
*+ bl_0_68 br_0_68 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c68
*+ bl_0_68 br_0_68 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c68
*+ bl_0_68 br_0_68 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c68
*+ bl_0_68 br_0_68 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c68
*+ bl_0_68 br_0_68 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c68
*+ bl_0_68 br_0_68 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c68
*+ bl_0_68 br_0_68 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c68
*+ bl_0_68 br_0_68 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c68
*+ bl_0_68 br_0_68 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c68
*+ bl_0_68 br_0_68 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c68
*+ bl_0_68 br_0_68 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c68
*+ bl_0_68 br_0_68 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c68
*+ bl_0_68 br_0_68 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c68
*+ bl_0_68 br_0_68 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c68
*+ bl_0_68 br_0_68 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c68
*+ bl_0_68 br_0_68 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c68
*+ bl_0_68 br_0_68 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c68
*+ bl_0_68 br_0_68 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c68
*+ bl_0_68 br_0_68 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c68
*+ bl_0_68 br_0_68 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c68
*+ bl_0_68 br_0_68 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c68
*+ bl_0_68 br_0_68 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c68
*+ bl_0_68 br_0_68 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c68
*+ bl_0_68 br_0_68 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c68
*+ bl_0_68 br_0_68 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c68
*+ bl_0_68 br_0_68 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c68
*+ bl_0_68 br_0_68 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c68
*+ bl_0_68 br_0_68 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c68
*+ bl_0_68 br_0_68 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c68
*+ bl_0_68 br_0_68 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c68
*+ bl_0_68 br_0_68 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c68
*+ bl_0_68 br_0_68 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c68
*+ bl_0_68 br_0_68 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c68
*+ bl_0_68 br_0_68 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c68
*+ bl_0_68 br_0_68 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c68
*+ bl_0_68 br_0_68 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c68
*+ bl_0_68 br_0_68 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c68
*+ bl_0_68 br_0_68 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c68
*+ bl_0_68 br_0_68 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c68
*+ bl_0_68 br_0_68 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c68
*+ bl_0_68 br_0_68 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c68
*+ bl_0_68 br_0_68 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c68
*+ bl_0_68 br_0_68 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c68
*+ bl_0_68 br_0_68 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c68
*+ bl_0_68 br_0_68 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c68
*+ bl_0_68 br_0_68 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c68
*+ bl_0_68 br_0_68 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c68
*+ bl_0_68 br_0_68 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c68
*+ bl_0_68 br_0_68 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c68
*+ bl_0_68 br_0_68 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c68
*+ bl_0_68 br_0_68 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c68
*+ bl_0_68 br_0_68 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c68
*+ bl_0_68 br_0_68 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c68
*+ bl_0_68 br_0_68 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c68
*+ bl_0_68 br_0_68 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c68
*+ bl_0_68 br_0_68 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c68
*+ bl_0_68 br_0_68 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c68
*+ bl_0_68 br_0_68 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c68
*+ bl_0_68 br_0_68 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c68
*+ bl_0_68 br_0_68 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c68
*+ bl_0_68 br_0_68 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c68
*+ bl_0_68 br_0_68 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c68
*+ bl_0_68 br_0_68 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c68
*+ bl_0_68 br_0_68 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c68
*+ bl_0_68 br_0_68 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c68
*+ bl_0_68 br_0_68 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c68
*+ bl_0_68 br_0_68 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c68
*+ bl_0_68 br_0_68 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c68
*+ bl_0_68 br_0_68 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c68
*+ bl_0_68 br_0_68 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c68
*+ bl_0_68 br_0_68 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c68
*+ bl_0_68 br_0_68 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c68
*+ bl_0_68 br_0_68 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c68
*+ bl_0_68 br_0_68 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c68
*+ bl_0_68 br_0_68 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c68
*+ bl_0_68 br_0_68 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c68
*+ bl_0_68 br_0_68 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c68
*+ bl_0_68 br_0_68 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c68
*+ bl_0_68 br_0_68 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c68
*+ bl_0_68 br_0_68 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c68
*+ bl_0_68 br_0_68 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c68
*+ bl_0_68 br_0_68 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c68
*+ bl_0_68 br_0_68 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c68
*+ bl_0_68 br_0_68 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c68
*+ bl_0_68 br_0_68 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c68
*+ bl_0_68 br_0_68 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c68
*+ bl_0_68 br_0_68 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c68
*+ bl_0_68 br_0_68 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c68
*+ bl_0_68 br_0_68 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c68
*+ bl_0_68 br_0_68 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c68
*+ bl_0_68 br_0_68 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c68
*+ bl_0_68 br_0_68 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c68
*+ bl_0_68 br_0_68 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c68
*+ bl_0_68 br_0_68 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c68
*+ bl_0_68 br_0_68 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c68
*+ bl_0_68 br_0_68 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c68
*+ bl_0_68 br_0_68 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c68
*+ bl_0_68 br_0_68 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c68
*+ bl_0_68 br_0_68 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c68
*+ bl_0_68 br_0_68 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c68
*+ bl_0_68 br_0_68 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c68
*+ bl_0_68 br_0_68 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c68
*+ bl_0_68 br_0_68 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c68
*+ bl_0_68 br_0_68 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c68
*+ bl_0_68 br_0_68 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c68
*+ bl_0_68 br_0_68 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c68
+ bl_0_68 br_0_68 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c69
+ bl_0_69 br_0_69 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c69
*+ bl_0_69 br_0_69 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c69
*+ bl_0_69 br_0_69 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c69
*+ bl_0_69 br_0_69 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c69
*+ bl_0_69 br_0_69 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c69
*+ bl_0_69 br_0_69 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c69
*+ bl_0_69 br_0_69 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c69
*+ bl_0_69 br_0_69 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c69
*+ bl_0_69 br_0_69 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c69
*+ bl_0_69 br_0_69 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c69
*+ bl_0_69 br_0_69 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c69
*+ bl_0_69 br_0_69 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c69
*+ bl_0_69 br_0_69 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c69
*+ bl_0_69 br_0_69 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c69
*+ bl_0_69 br_0_69 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c69
*+ bl_0_69 br_0_69 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c69
*+ bl_0_69 br_0_69 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c69
*+ bl_0_69 br_0_69 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c69
*+ bl_0_69 br_0_69 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c69
*+ bl_0_69 br_0_69 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c69
*+ bl_0_69 br_0_69 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c69
*+ bl_0_69 br_0_69 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c69
*+ bl_0_69 br_0_69 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c69
*+ bl_0_69 br_0_69 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c69
*+ bl_0_69 br_0_69 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c69
*+ bl_0_69 br_0_69 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c69
*+ bl_0_69 br_0_69 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c69
*+ bl_0_69 br_0_69 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c69
*+ bl_0_69 br_0_69 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c69
*+ bl_0_69 br_0_69 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c69
*+ bl_0_69 br_0_69 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c69
*+ bl_0_69 br_0_69 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c69
*+ bl_0_69 br_0_69 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c69
*+ bl_0_69 br_0_69 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c69
*+ bl_0_69 br_0_69 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c69
*+ bl_0_69 br_0_69 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c69
*+ bl_0_69 br_0_69 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c69
*+ bl_0_69 br_0_69 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c69
*+ bl_0_69 br_0_69 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c69
*+ bl_0_69 br_0_69 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c69
*+ bl_0_69 br_0_69 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c69
*+ bl_0_69 br_0_69 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c69
*+ bl_0_69 br_0_69 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c69
*+ bl_0_69 br_0_69 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c69
*+ bl_0_69 br_0_69 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c69
*+ bl_0_69 br_0_69 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c69
*+ bl_0_69 br_0_69 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c69
*+ bl_0_69 br_0_69 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c69
*+ bl_0_69 br_0_69 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c69
*+ bl_0_69 br_0_69 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c69
*+ bl_0_69 br_0_69 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c69
*+ bl_0_69 br_0_69 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c69
*+ bl_0_69 br_0_69 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c69
*+ bl_0_69 br_0_69 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c69
*+ bl_0_69 br_0_69 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c69
*+ bl_0_69 br_0_69 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c69
*+ bl_0_69 br_0_69 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c69
*+ bl_0_69 br_0_69 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c69
*+ bl_0_69 br_0_69 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c69
*+ bl_0_69 br_0_69 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c69
*+ bl_0_69 br_0_69 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c69
*+ bl_0_69 br_0_69 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c69
*+ bl_0_69 br_0_69 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c69
*+ bl_0_69 br_0_69 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c69
*+ bl_0_69 br_0_69 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c69
*+ bl_0_69 br_0_69 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c69
*+ bl_0_69 br_0_69 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c69
*+ bl_0_69 br_0_69 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c69
*+ bl_0_69 br_0_69 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c69
*+ bl_0_69 br_0_69 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c69
*+ bl_0_69 br_0_69 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c69
*+ bl_0_69 br_0_69 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c69
*+ bl_0_69 br_0_69 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c69
*+ bl_0_69 br_0_69 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c69
*+ bl_0_69 br_0_69 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c69
*+ bl_0_69 br_0_69 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c69
*+ bl_0_69 br_0_69 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c69
*+ bl_0_69 br_0_69 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c69
*+ bl_0_69 br_0_69 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c69
*+ bl_0_69 br_0_69 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c69
*+ bl_0_69 br_0_69 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c69
*+ bl_0_69 br_0_69 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c69
*+ bl_0_69 br_0_69 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c69
*+ bl_0_69 br_0_69 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c69
*+ bl_0_69 br_0_69 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c69
*+ bl_0_69 br_0_69 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c69
*+ bl_0_69 br_0_69 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c69
*+ bl_0_69 br_0_69 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c69
*+ bl_0_69 br_0_69 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c69
*+ bl_0_69 br_0_69 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c69
*+ bl_0_69 br_0_69 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c69
*+ bl_0_69 br_0_69 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c69
*+ bl_0_69 br_0_69 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c69
*+ bl_0_69 br_0_69 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c69
*+ bl_0_69 br_0_69 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c69
*+ bl_0_69 br_0_69 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c69
*+ bl_0_69 br_0_69 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c69
*+ bl_0_69 br_0_69 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c69
*+ bl_0_69 br_0_69 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c69
*+ bl_0_69 br_0_69 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c69
*+ bl_0_69 br_0_69 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c69
*+ bl_0_69 br_0_69 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c69
*+ bl_0_69 br_0_69 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c69
*+ bl_0_69 br_0_69 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c69
*+ bl_0_69 br_0_69 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c69
*+ bl_0_69 br_0_69 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c69
*+ bl_0_69 br_0_69 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c69
*+ bl_0_69 br_0_69 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c69
*+ bl_0_69 br_0_69 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c69
*+ bl_0_69 br_0_69 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c69
*+ bl_0_69 br_0_69 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c69
*+ bl_0_69 br_0_69 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c69
*+ bl_0_69 br_0_69 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c69
*+ bl_0_69 br_0_69 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c69
*+ bl_0_69 br_0_69 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c69
*+ bl_0_69 br_0_69 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c69
*+ bl_0_69 br_0_69 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c69
*+ bl_0_69 br_0_69 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c69
*+ bl_0_69 br_0_69 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c69
*+ bl_0_69 br_0_69 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c69
*+ bl_0_69 br_0_69 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c69
*+ bl_0_69 br_0_69 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c69
*+ bl_0_69 br_0_69 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c69
*+ bl_0_69 br_0_69 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c69
*+ bl_0_69 br_0_69 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c69
*+ bl_0_69 br_0_69 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c69
*+ bl_0_69 br_0_69 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c69
+ bl_0_69 br_0_69 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c70
+ bl_0_70 br_0_70 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c70
*+ bl_0_70 br_0_70 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c70
*+ bl_0_70 br_0_70 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c70
*+ bl_0_70 br_0_70 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c70
*+ bl_0_70 br_0_70 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c70
*+ bl_0_70 br_0_70 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c70
*+ bl_0_70 br_0_70 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c70
*+ bl_0_70 br_0_70 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c70
*+ bl_0_70 br_0_70 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c70
*+ bl_0_70 br_0_70 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c70
*+ bl_0_70 br_0_70 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c70
*+ bl_0_70 br_0_70 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c70
*+ bl_0_70 br_0_70 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c70
*+ bl_0_70 br_0_70 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c70
*+ bl_0_70 br_0_70 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c70
*+ bl_0_70 br_0_70 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c70
*+ bl_0_70 br_0_70 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c70
*+ bl_0_70 br_0_70 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c70
*+ bl_0_70 br_0_70 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c70
*+ bl_0_70 br_0_70 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c70
*+ bl_0_70 br_0_70 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c70
*+ bl_0_70 br_0_70 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c70
*+ bl_0_70 br_0_70 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c70
*+ bl_0_70 br_0_70 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c70
*+ bl_0_70 br_0_70 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c70
*+ bl_0_70 br_0_70 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c70
*+ bl_0_70 br_0_70 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c70
*+ bl_0_70 br_0_70 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c70
*+ bl_0_70 br_0_70 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c70
*+ bl_0_70 br_0_70 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c70
*+ bl_0_70 br_0_70 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c70
*+ bl_0_70 br_0_70 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c70
*+ bl_0_70 br_0_70 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c70
*+ bl_0_70 br_0_70 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c70
*+ bl_0_70 br_0_70 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c70
*+ bl_0_70 br_0_70 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c70
*+ bl_0_70 br_0_70 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c70
*+ bl_0_70 br_0_70 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c70
*+ bl_0_70 br_0_70 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c70
*+ bl_0_70 br_0_70 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c70
*+ bl_0_70 br_0_70 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c70
*+ bl_0_70 br_0_70 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c70
*+ bl_0_70 br_0_70 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c70
*+ bl_0_70 br_0_70 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c70
*+ bl_0_70 br_0_70 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c70
*+ bl_0_70 br_0_70 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c70
*+ bl_0_70 br_0_70 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c70
*+ bl_0_70 br_0_70 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c70
*+ bl_0_70 br_0_70 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c70
*+ bl_0_70 br_0_70 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c70
*+ bl_0_70 br_0_70 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c70
*+ bl_0_70 br_0_70 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c70
*+ bl_0_70 br_0_70 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c70
*+ bl_0_70 br_0_70 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c70
*+ bl_0_70 br_0_70 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c70
*+ bl_0_70 br_0_70 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c70
*+ bl_0_70 br_0_70 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c70
*+ bl_0_70 br_0_70 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c70
*+ bl_0_70 br_0_70 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c70
*+ bl_0_70 br_0_70 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c70
*+ bl_0_70 br_0_70 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c70
*+ bl_0_70 br_0_70 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c70
*+ bl_0_70 br_0_70 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c70
*+ bl_0_70 br_0_70 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c70
*+ bl_0_70 br_0_70 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c70
*+ bl_0_70 br_0_70 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c70
*+ bl_0_70 br_0_70 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c70
*+ bl_0_70 br_0_70 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c70
*+ bl_0_70 br_0_70 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c70
*+ bl_0_70 br_0_70 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c70
*+ bl_0_70 br_0_70 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c70
*+ bl_0_70 br_0_70 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c70
*+ bl_0_70 br_0_70 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c70
*+ bl_0_70 br_0_70 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c70
*+ bl_0_70 br_0_70 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c70
*+ bl_0_70 br_0_70 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c70
*+ bl_0_70 br_0_70 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c70
*+ bl_0_70 br_0_70 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c70
*+ bl_0_70 br_0_70 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c70
*+ bl_0_70 br_0_70 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c70
*+ bl_0_70 br_0_70 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c70
*+ bl_0_70 br_0_70 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c70
*+ bl_0_70 br_0_70 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c70
*+ bl_0_70 br_0_70 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c70
*+ bl_0_70 br_0_70 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c70
*+ bl_0_70 br_0_70 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c70
*+ bl_0_70 br_0_70 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c70
*+ bl_0_70 br_0_70 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c70
*+ bl_0_70 br_0_70 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c70
*+ bl_0_70 br_0_70 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c70
*+ bl_0_70 br_0_70 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c70
*+ bl_0_70 br_0_70 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c70
*+ bl_0_70 br_0_70 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c70
*+ bl_0_70 br_0_70 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c70
*+ bl_0_70 br_0_70 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c70
*+ bl_0_70 br_0_70 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c70
*+ bl_0_70 br_0_70 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c70
*+ bl_0_70 br_0_70 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c70
*+ bl_0_70 br_0_70 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c70
*+ bl_0_70 br_0_70 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c70
*+ bl_0_70 br_0_70 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c70
*+ bl_0_70 br_0_70 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c70
*+ bl_0_70 br_0_70 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c70
*+ bl_0_70 br_0_70 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c70
*+ bl_0_70 br_0_70 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c70
*+ bl_0_70 br_0_70 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c70
*+ bl_0_70 br_0_70 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c70
*+ bl_0_70 br_0_70 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c70
*+ bl_0_70 br_0_70 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c70
*+ bl_0_70 br_0_70 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c70
*+ bl_0_70 br_0_70 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c70
*+ bl_0_70 br_0_70 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c70
*+ bl_0_70 br_0_70 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c70
*+ bl_0_70 br_0_70 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c70
*+ bl_0_70 br_0_70 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c70
*+ bl_0_70 br_0_70 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c70
*+ bl_0_70 br_0_70 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c70
*+ bl_0_70 br_0_70 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c70
*+ bl_0_70 br_0_70 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c70
*+ bl_0_70 br_0_70 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c70
*+ bl_0_70 br_0_70 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c70
*+ bl_0_70 br_0_70 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c70
*+ bl_0_70 br_0_70 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c70
*+ bl_0_70 br_0_70 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c70
*+ bl_0_70 br_0_70 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c70
*+ bl_0_70 br_0_70 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c70
*+ bl_0_70 br_0_70 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c70
+ bl_0_70 br_0_70 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c71
+ bl_0_71 br_0_71 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c71
*+ bl_0_71 br_0_71 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c71
*+ bl_0_71 br_0_71 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c71
*+ bl_0_71 br_0_71 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c71
*+ bl_0_71 br_0_71 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c71
*+ bl_0_71 br_0_71 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c71
*+ bl_0_71 br_0_71 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c71
*+ bl_0_71 br_0_71 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c71
*+ bl_0_71 br_0_71 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c71
*+ bl_0_71 br_0_71 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c71
*+ bl_0_71 br_0_71 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c71
*+ bl_0_71 br_0_71 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c71
*+ bl_0_71 br_0_71 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c71
*+ bl_0_71 br_0_71 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c71
*+ bl_0_71 br_0_71 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c71
*+ bl_0_71 br_0_71 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c71
*+ bl_0_71 br_0_71 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c71
*+ bl_0_71 br_0_71 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c71
*+ bl_0_71 br_0_71 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c71
*+ bl_0_71 br_0_71 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c71
*+ bl_0_71 br_0_71 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c71
*+ bl_0_71 br_0_71 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c71
*+ bl_0_71 br_0_71 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c71
*+ bl_0_71 br_0_71 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c71
*+ bl_0_71 br_0_71 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c71
*+ bl_0_71 br_0_71 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c71
*+ bl_0_71 br_0_71 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c71
*+ bl_0_71 br_0_71 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c71
*+ bl_0_71 br_0_71 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c71
*+ bl_0_71 br_0_71 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c71
*+ bl_0_71 br_0_71 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c71
*+ bl_0_71 br_0_71 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c71
*+ bl_0_71 br_0_71 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c71
*+ bl_0_71 br_0_71 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c71
*+ bl_0_71 br_0_71 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c71
*+ bl_0_71 br_0_71 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c71
*+ bl_0_71 br_0_71 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c71
*+ bl_0_71 br_0_71 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c71
*+ bl_0_71 br_0_71 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c71
*+ bl_0_71 br_0_71 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c71
*+ bl_0_71 br_0_71 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c71
*+ bl_0_71 br_0_71 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c71
*+ bl_0_71 br_0_71 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c71
*+ bl_0_71 br_0_71 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c71
*+ bl_0_71 br_0_71 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c71
*+ bl_0_71 br_0_71 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c71
*+ bl_0_71 br_0_71 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c71
*+ bl_0_71 br_0_71 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c71
*+ bl_0_71 br_0_71 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c71
*+ bl_0_71 br_0_71 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c71
*+ bl_0_71 br_0_71 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c71
*+ bl_0_71 br_0_71 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c71
*+ bl_0_71 br_0_71 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c71
*+ bl_0_71 br_0_71 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c71
*+ bl_0_71 br_0_71 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c71
*+ bl_0_71 br_0_71 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c71
*+ bl_0_71 br_0_71 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c71
*+ bl_0_71 br_0_71 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c71
*+ bl_0_71 br_0_71 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c71
*+ bl_0_71 br_0_71 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c71
*+ bl_0_71 br_0_71 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c71
*+ bl_0_71 br_0_71 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c71
*+ bl_0_71 br_0_71 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c71
*+ bl_0_71 br_0_71 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c71
*+ bl_0_71 br_0_71 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c71
*+ bl_0_71 br_0_71 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c71
*+ bl_0_71 br_0_71 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c71
*+ bl_0_71 br_0_71 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c71
*+ bl_0_71 br_0_71 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c71
*+ bl_0_71 br_0_71 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c71
*+ bl_0_71 br_0_71 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c71
*+ bl_0_71 br_0_71 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c71
*+ bl_0_71 br_0_71 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c71
*+ bl_0_71 br_0_71 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c71
*+ bl_0_71 br_0_71 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c71
*+ bl_0_71 br_0_71 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c71
*+ bl_0_71 br_0_71 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c71
*+ bl_0_71 br_0_71 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c71
*+ bl_0_71 br_0_71 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c71
*+ bl_0_71 br_0_71 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c71
*+ bl_0_71 br_0_71 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c71
*+ bl_0_71 br_0_71 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c71
*+ bl_0_71 br_0_71 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c71
*+ bl_0_71 br_0_71 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c71
*+ bl_0_71 br_0_71 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c71
*+ bl_0_71 br_0_71 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c71
*+ bl_0_71 br_0_71 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c71
*+ bl_0_71 br_0_71 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c71
*+ bl_0_71 br_0_71 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c71
*+ bl_0_71 br_0_71 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c71
*+ bl_0_71 br_0_71 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c71
*+ bl_0_71 br_0_71 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c71
*+ bl_0_71 br_0_71 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c71
*+ bl_0_71 br_0_71 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c71
*+ bl_0_71 br_0_71 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c71
*+ bl_0_71 br_0_71 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c71
*+ bl_0_71 br_0_71 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c71
*+ bl_0_71 br_0_71 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c71
*+ bl_0_71 br_0_71 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c71
*+ bl_0_71 br_0_71 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c71
*+ bl_0_71 br_0_71 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c71
*+ bl_0_71 br_0_71 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c71
*+ bl_0_71 br_0_71 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c71
*+ bl_0_71 br_0_71 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c71
*+ bl_0_71 br_0_71 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c71
*+ bl_0_71 br_0_71 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c71
*+ bl_0_71 br_0_71 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c71
*+ bl_0_71 br_0_71 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c71
*+ bl_0_71 br_0_71 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c71
*+ bl_0_71 br_0_71 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c71
*+ bl_0_71 br_0_71 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c71
*+ bl_0_71 br_0_71 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c71
*+ bl_0_71 br_0_71 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c71
*+ bl_0_71 br_0_71 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c71
*+ bl_0_71 br_0_71 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c71
*+ bl_0_71 br_0_71 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c71
*+ bl_0_71 br_0_71 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c71
*+ bl_0_71 br_0_71 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c71
*+ bl_0_71 br_0_71 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c71
*+ bl_0_71 br_0_71 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c71
*+ bl_0_71 br_0_71 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c71
*+ bl_0_71 br_0_71 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c71
*+ bl_0_71 br_0_71 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c71
*+ bl_0_71 br_0_71 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c71
*+ bl_0_71 br_0_71 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c71
*+ bl_0_71 br_0_71 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c71
*+ bl_0_71 br_0_71 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c71
+ bl_0_71 br_0_71 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c72
+ bl_0_72 br_0_72 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c72
*+ bl_0_72 br_0_72 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c72
*+ bl_0_72 br_0_72 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c72
*+ bl_0_72 br_0_72 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c72
*+ bl_0_72 br_0_72 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c72
*+ bl_0_72 br_0_72 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c72
*+ bl_0_72 br_0_72 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c72
*+ bl_0_72 br_0_72 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c72
*+ bl_0_72 br_0_72 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c72
*+ bl_0_72 br_0_72 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c72
*+ bl_0_72 br_0_72 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c72
*+ bl_0_72 br_0_72 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c72
*+ bl_0_72 br_0_72 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c72
*+ bl_0_72 br_0_72 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c72
*+ bl_0_72 br_0_72 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c72
*+ bl_0_72 br_0_72 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c72
*+ bl_0_72 br_0_72 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c72
*+ bl_0_72 br_0_72 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c72
*+ bl_0_72 br_0_72 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c72
*+ bl_0_72 br_0_72 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c72
*+ bl_0_72 br_0_72 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c72
*+ bl_0_72 br_0_72 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c72
*+ bl_0_72 br_0_72 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c72
*+ bl_0_72 br_0_72 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c72
*+ bl_0_72 br_0_72 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c72
*+ bl_0_72 br_0_72 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c72
*+ bl_0_72 br_0_72 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c72
*+ bl_0_72 br_0_72 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c72
*+ bl_0_72 br_0_72 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c72
*+ bl_0_72 br_0_72 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c72
*+ bl_0_72 br_0_72 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c72
*+ bl_0_72 br_0_72 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c72
*+ bl_0_72 br_0_72 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c72
*+ bl_0_72 br_0_72 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c72
*+ bl_0_72 br_0_72 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c72
*+ bl_0_72 br_0_72 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c72
*+ bl_0_72 br_0_72 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c72
*+ bl_0_72 br_0_72 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c72
*+ bl_0_72 br_0_72 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c72
*+ bl_0_72 br_0_72 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c72
*+ bl_0_72 br_0_72 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c72
*+ bl_0_72 br_0_72 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c72
*+ bl_0_72 br_0_72 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c72
*+ bl_0_72 br_0_72 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c72
*+ bl_0_72 br_0_72 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c72
*+ bl_0_72 br_0_72 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c72
*+ bl_0_72 br_0_72 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c72
*+ bl_0_72 br_0_72 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c72
*+ bl_0_72 br_0_72 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c72
*+ bl_0_72 br_0_72 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c72
*+ bl_0_72 br_0_72 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c72
*+ bl_0_72 br_0_72 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c72
*+ bl_0_72 br_0_72 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c72
*+ bl_0_72 br_0_72 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c72
*+ bl_0_72 br_0_72 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c72
*+ bl_0_72 br_0_72 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c72
*+ bl_0_72 br_0_72 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c72
*+ bl_0_72 br_0_72 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c72
*+ bl_0_72 br_0_72 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c72
*+ bl_0_72 br_0_72 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c72
*+ bl_0_72 br_0_72 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c72
*+ bl_0_72 br_0_72 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c72
*+ bl_0_72 br_0_72 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c72
*+ bl_0_72 br_0_72 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c72
*+ bl_0_72 br_0_72 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c72
*+ bl_0_72 br_0_72 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c72
*+ bl_0_72 br_0_72 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c72
*+ bl_0_72 br_0_72 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c72
*+ bl_0_72 br_0_72 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c72
*+ bl_0_72 br_0_72 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c72
*+ bl_0_72 br_0_72 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c72
*+ bl_0_72 br_0_72 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c72
*+ bl_0_72 br_0_72 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c72
*+ bl_0_72 br_0_72 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c72
*+ bl_0_72 br_0_72 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c72
*+ bl_0_72 br_0_72 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c72
*+ bl_0_72 br_0_72 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c72
*+ bl_0_72 br_0_72 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c72
*+ bl_0_72 br_0_72 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c72
*+ bl_0_72 br_0_72 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c72
*+ bl_0_72 br_0_72 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c72
*+ bl_0_72 br_0_72 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c72
*+ bl_0_72 br_0_72 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c72
*+ bl_0_72 br_0_72 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c72
*+ bl_0_72 br_0_72 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c72
*+ bl_0_72 br_0_72 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c72
*+ bl_0_72 br_0_72 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c72
*+ bl_0_72 br_0_72 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c72
*+ bl_0_72 br_0_72 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c72
*+ bl_0_72 br_0_72 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c72
*+ bl_0_72 br_0_72 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c72
*+ bl_0_72 br_0_72 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c72
*+ bl_0_72 br_0_72 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c72
*+ bl_0_72 br_0_72 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c72
*+ bl_0_72 br_0_72 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c72
*+ bl_0_72 br_0_72 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c72
*+ bl_0_72 br_0_72 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c72
*+ bl_0_72 br_0_72 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c72
*+ bl_0_72 br_0_72 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c72
*+ bl_0_72 br_0_72 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c72
*+ bl_0_72 br_0_72 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c72
*+ bl_0_72 br_0_72 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c72
*+ bl_0_72 br_0_72 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c72
*+ bl_0_72 br_0_72 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c72
*+ bl_0_72 br_0_72 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c72
*+ bl_0_72 br_0_72 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c72
*+ bl_0_72 br_0_72 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c72
*+ bl_0_72 br_0_72 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c72
*+ bl_0_72 br_0_72 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c72
*+ bl_0_72 br_0_72 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c72
*+ bl_0_72 br_0_72 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c72
*+ bl_0_72 br_0_72 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c72
*+ bl_0_72 br_0_72 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c72
*+ bl_0_72 br_0_72 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c72
*+ bl_0_72 br_0_72 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c72
*+ bl_0_72 br_0_72 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c72
*+ bl_0_72 br_0_72 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c72
*+ bl_0_72 br_0_72 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c72
*+ bl_0_72 br_0_72 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c72
*+ bl_0_72 br_0_72 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c72
*+ bl_0_72 br_0_72 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c72
*+ bl_0_72 br_0_72 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c72
*+ bl_0_72 br_0_72 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c72
*+ bl_0_72 br_0_72 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c72
*+ bl_0_72 br_0_72 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c72
*+ bl_0_72 br_0_72 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c72
*+ bl_0_72 br_0_72 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c72
+ bl_0_72 br_0_72 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c73
+ bl_0_73 br_0_73 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c73
*+ bl_0_73 br_0_73 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c73
*+ bl_0_73 br_0_73 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c73
*+ bl_0_73 br_0_73 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c73
*+ bl_0_73 br_0_73 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c73
*+ bl_0_73 br_0_73 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c73
*+ bl_0_73 br_0_73 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c73
*+ bl_0_73 br_0_73 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c73
*+ bl_0_73 br_0_73 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c73
*+ bl_0_73 br_0_73 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c73
*+ bl_0_73 br_0_73 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c73
*+ bl_0_73 br_0_73 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c73
*+ bl_0_73 br_0_73 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c73
*+ bl_0_73 br_0_73 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c73
*+ bl_0_73 br_0_73 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c73
*+ bl_0_73 br_0_73 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c73
*+ bl_0_73 br_0_73 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c73
*+ bl_0_73 br_0_73 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c73
*+ bl_0_73 br_0_73 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c73
*+ bl_0_73 br_0_73 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c73
*+ bl_0_73 br_0_73 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c73
*+ bl_0_73 br_0_73 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c73
*+ bl_0_73 br_0_73 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c73
*+ bl_0_73 br_0_73 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c73
*+ bl_0_73 br_0_73 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c73
*+ bl_0_73 br_0_73 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c73
*+ bl_0_73 br_0_73 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c73
*+ bl_0_73 br_0_73 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c73
*+ bl_0_73 br_0_73 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c73
*+ bl_0_73 br_0_73 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c73
*+ bl_0_73 br_0_73 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c73
*+ bl_0_73 br_0_73 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c73
*+ bl_0_73 br_0_73 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c73
*+ bl_0_73 br_0_73 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c73
*+ bl_0_73 br_0_73 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c73
*+ bl_0_73 br_0_73 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c73
*+ bl_0_73 br_0_73 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c73
*+ bl_0_73 br_0_73 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c73
*+ bl_0_73 br_0_73 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c73
*+ bl_0_73 br_0_73 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c73
*+ bl_0_73 br_0_73 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c73
*+ bl_0_73 br_0_73 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c73
*+ bl_0_73 br_0_73 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c73
*+ bl_0_73 br_0_73 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c73
*+ bl_0_73 br_0_73 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c73
*+ bl_0_73 br_0_73 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c73
*+ bl_0_73 br_0_73 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c73
*+ bl_0_73 br_0_73 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c73
*+ bl_0_73 br_0_73 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c73
*+ bl_0_73 br_0_73 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c73
*+ bl_0_73 br_0_73 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c73
*+ bl_0_73 br_0_73 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c73
*+ bl_0_73 br_0_73 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c73
*+ bl_0_73 br_0_73 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c73
*+ bl_0_73 br_0_73 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c73
*+ bl_0_73 br_0_73 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c73
*+ bl_0_73 br_0_73 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c73
*+ bl_0_73 br_0_73 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c73
*+ bl_0_73 br_0_73 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c73
*+ bl_0_73 br_0_73 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c73
*+ bl_0_73 br_0_73 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c73
*+ bl_0_73 br_0_73 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c73
*+ bl_0_73 br_0_73 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c73
*+ bl_0_73 br_0_73 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c73
*+ bl_0_73 br_0_73 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c73
*+ bl_0_73 br_0_73 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c73
*+ bl_0_73 br_0_73 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c73
*+ bl_0_73 br_0_73 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c73
*+ bl_0_73 br_0_73 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c73
*+ bl_0_73 br_0_73 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c73
*+ bl_0_73 br_0_73 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c73
*+ bl_0_73 br_0_73 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c73
*+ bl_0_73 br_0_73 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c73
*+ bl_0_73 br_0_73 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c73
*+ bl_0_73 br_0_73 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c73
*+ bl_0_73 br_0_73 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c73
*+ bl_0_73 br_0_73 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c73
*+ bl_0_73 br_0_73 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c73
*+ bl_0_73 br_0_73 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c73
*+ bl_0_73 br_0_73 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c73
*+ bl_0_73 br_0_73 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c73
*+ bl_0_73 br_0_73 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c73
*+ bl_0_73 br_0_73 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c73
*+ bl_0_73 br_0_73 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c73
*+ bl_0_73 br_0_73 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c73
*+ bl_0_73 br_0_73 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c73
*+ bl_0_73 br_0_73 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c73
*+ bl_0_73 br_0_73 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c73
*+ bl_0_73 br_0_73 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c73
*+ bl_0_73 br_0_73 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c73
*+ bl_0_73 br_0_73 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c73
*+ bl_0_73 br_0_73 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c73
*+ bl_0_73 br_0_73 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c73
*+ bl_0_73 br_0_73 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c73
*+ bl_0_73 br_0_73 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c73
*+ bl_0_73 br_0_73 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c73
*+ bl_0_73 br_0_73 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c73
*+ bl_0_73 br_0_73 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c73
*+ bl_0_73 br_0_73 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c73
*+ bl_0_73 br_0_73 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c73
*+ bl_0_73 br_0_73 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c73
*+ bl_0_73 br_0_73 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c73
*+ bl_0_73 br_0_73 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c73
*+ bl_0_73 br_0_73 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c73
*+ bl_0_73 br_0_73 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c73
*+ bl_0_73 br_0_73 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c73
*+ bl_0_73 br_0_73 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c73
*+ bl_0_73 br_0_73 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c73
*+ bl_0_73 br_0_73 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c73
*+ bl_0_73 br_0_73 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c73
*+ bl_0_73 br_0_73 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c73
*+ bl_0_73 br_0_73 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c73
*+ bl_0_73 br_0_73 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c73
*+ bl_0_73 br_0_73 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c73
*+ bl_0_73 br_0_73 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c73
*+ bl_0_73 br_0_73 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c73
*+ bl_0_73 br_0_73 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c73
*+ bl_0_73 br_0_73 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c73
*+ bl_0_73 br_0_73 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c73
*+ bl_0_73 br_0_73 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c73
*+ bl_0_73 br_0_73 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c73
*+ bl_0_73 br_0_73 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c73
*+ bl_0_73 br_0_73 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c73
*+ bl_0_73 br_0_73 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c73
*+ bl_0_73 br_0_73 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c73
*+ bl_0_73 br_0_73 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c73
*+ bl_0_73 br_0_73 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c73
+ bl_0_73 br_0_73 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c74
+ bl_0_74 br_0_74 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c74
*+ bl_0_74 br_0_74 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c74
*+ bl_0_74 br_0_74 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c74
*+ bl_0_74 br_0_74 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c74
*+ bl_0_74 br_0_74 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c74
*+ bl_0_74 br_0_74 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c74
*+ bl_0_74 br_0_74 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c74
*+ bl_0_74 br_0_74 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c74
*+ bl_0_74 br_0_74 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c74
*+ bl_0_74 br_0_74 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c74
*+ bl_0_74 br_0_74 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c74
*+ bl_0_74 br_0_74 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c74
*+ bl_0_74 br_0_74 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c74
*+ bl_0_74 br_0_74 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c74
*+ bl_0_74 br_0_74 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c74
*+ bl_0_74 br_0_74 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c74
*+ bl_0_74 br_0_74 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c74
*+ bl_0_74 br_0_74 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c74
*+ bl_0_74 br_0_74 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c74
*+ bl_0_74 br_0_74 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c74
*+ bl_0_74 br_0_74 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c74
*+ bl_0_74 br_0_74 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c74
*+ bl_0_74 br_0_74 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c74
*+ bl_0_74 br_0_74 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c74
*+ bl_0_74 br_0_74 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c74
*+ bl_0_74 br_0_74 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c74
*+ bl_0_74 br_0_74 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c74
*+ bl_0_74 br_0_74 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c74
*+ bl_0_74 br_0_74 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c74
*+ bl_0_74 br_0_74 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c74
*+ bl_0_74 br_0_74 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c74
*+ bl_0_74 br_0_74 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c74
*+ bl_0_74 br_0_74 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c74
*+ bl_0_74 br_0_74 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c74
*+ bl_0_74 br_0_74 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c74
*+ bl_0_74 br_0_74 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c74
*+ bl_0_74 br_0_74 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c74
*+ bl_0_74 br_0_74 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c74
*+ bl_0_74 br_0_74 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c74
*+ bl_0_74 br_0_74 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c74
*+ bl_0_74 br_0_74 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c74
*+ bl_0_74 br_0_74 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c74
*+ bl_0_74 br_0_74 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c74
*+ bl_0_74 br_0_74 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c74
*+ bl_0_74 br_0_74 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c74
*+ bl_0_74 br_0_74 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c74
*+ bl_0_74 br_0_74 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c74
*+ bl_0_74 br_0_74 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c74
*+ bl_0_74 br_0_74 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c74
*+ bl_0_74 br_0_74 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c74
*+ bl_0_74 br_0_74 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c74
*+ bl_0_74 br_0_74 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c74
*+ bl_0_74 br_0_74 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c74
*+ bl_0_74 br_0_74 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c74
*+ bl_0_74 br_0_74 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c74
*+ bl_0_74 br_0_74 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c74
*+ bl_0_74 br_0_74 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c74
*+ bl_0_74 br_0_74 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c74
*+ bl_0_74 br_0_74 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c74
*+ bl_0_74 br_0_74 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c74
*+ bl_0_74 br_0_74 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c74
*+ bl_0_74 br_0_74 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c74
*+ bl_0_74 br_0_74 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c74
*+ bl_0_74 br_0_74 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c74
*+ bl_0_74 br_0_74 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c74
*+ bl_0_74 br_0_74 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c74
*+ bl_0_74 br_0_74 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c74
*+ bl_0_74 br_0_74 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c74
*+ bl_0_74 br_0_74 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c74
*+ bl_0_74 br_0_74 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c74
*+ bl_0_74 br_0_74 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c74
*+ bl_0_74 br_0_74 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c74
*+ bl_0_74 br_0_74 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c74
*+ bl_0_74 br_0_74 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c74
*+ bl_0_74 br_0_74 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c74
*+ bl_0_74 br_0_74 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c74
*+ bl_0_74 br_0_74 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c74
*+ bl_0_74 br_0_74 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c74
*+ bl_0_74 br_0_74 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c74
*+ bl_0_74 br_0_74 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c74
*+ bl_0_74 br_0_74 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c74
*+ bl_0_74 br_0_74 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c74
*+ bl_0_74 br_0_74 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c74
*+ bl_0_74 br_0_74 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c74
*+ bl_0_74 br_0_74 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c74
*+ bl_0_74 br_0_74 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c74
*+ bl_0_74 br_0_74 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c74
*+ bl_0_74 br_0_74 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c74
*+ bl_0_74 br_0_74 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c74
*+ bl_0_74 br_0_74 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c74
*+ bl_0_74 br_0_74 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c74
*+ bl_0_74 br_0_74 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c74
*+ bl_0_74 br_0_74 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c74
*+ bl_0_74 br_0_74 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c74
*+ bl_0_74 br_0_74 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c74
*+ bl_0_74 br_0_74 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c74
*+ bl_0_74 br_0_74 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c74
*+ bl_0_74 br_0_74 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c74
*+ bl_0_74 br_0_74 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c74
*+ bl_0_74 br_0_74 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c74
*+ bl_0_74 br_0_74 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c74
*+ bl_0_74 br_0_74 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c74
*+ bl_0_74 br_0_74 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c74
*+ bl_0_74 br_0_74 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c74
*+ bl_0_74 br_0_74 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c74
*+ bl_0_74 br_0_74 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c74
*+ bl_0_74 br_0_74 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c74
*+ bl_0_74 br_0_74 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c74
*+ bl_0_74 br_0_74 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c74
*+ bl_0_74 br_0_74 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c74
*+ bl_0_74 br_0_74 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c74
*+ bl_0_74 br_0_74 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c74
*+ bl_0_74 br_0_74 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c74
*+ bl_0_74 br_0_74 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c74
*+ bl_0_74 br_0_74 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c74
*+ bl_0_74 br_0_74 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c74
*+ bl_0_74 br_0_74 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c74
*+ bl_0_74 br_0_74 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c74
*+ bl_0_74 br_0_74 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c74
*+ bl_0_74 br_0_74 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c74
*+ bl_0_74 br_0_74 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c74
*+ bl_0_74 br_0_74 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c74
*+ bl_0_74 br_0_74 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c74
*+ bl_0_74 br_0_74 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c74
*+ bl_0_74 br_0_74 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c74
*+ bl_0_74 br_0_74 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c74
*+ bl_0_74 br_0_74 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c74
+ bl_0_74 br_0_74 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c75
+ bl_0_75 br_0_75 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c75
*+ bl_0_75 br_0_75 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c75
*+ bl_0_75 br_0_75 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c75
*+ bl_0_75 br_0_75 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c75
*+ bl_0_75 br_0_75 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c75
*+ bl_0_75 br_0_75 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c75
*+ bl_0_75 br_0_75 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c75
*+ bl_0_75 br_0_75 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c75
*+ bl_0_75 br_0_75 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c75
*+ bl_0_75 br_0_75 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c75
*+ bl_0_75 br_0_75 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c75
*+ bl_0_75 br_0_75 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c75
*+ bl_0_75 br_0_75 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c75
*+ bl_0_75 br_0_75 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c75
*+ bl_0_75 br_0_75 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c75
*+ bl_0_75 br_0_75 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c75
*+ bl_0_75 br_0_75 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c75
*+ bl_0_75 br_0_75 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c75
*+ bl_0_75 br_0_75 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c75
*+ bl_0_75 br_0_75 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c75
*+ bl_0_75 br_0_75 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c75
*+ bl_0_75 br_0_75 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c75
*+ bl_0_75 br_0_75 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c75
*+ bl_0_75 br_0_75 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c75
*+ bl_0_75 br_0_75 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c75
*+ bl_0_75 br_0_75 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c75
*+ bl_0_75 br_0_75 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c75
*+ bl_0_75 br_0_75 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c75
*+ bl_0_75 br_0_75 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c75
*+ bl_0_75 br_0_75 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c75
*+ bl_0_75 br_0_75 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c75
*+ bl_0_75 br_0_75 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c75
*+ bl_0_75 br_0_75 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c75
*+ bl_0_75 br_0_75 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c75
*+ bl_0_75 br_0_75 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c75
*+ bl_0_75 br_0_75 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c75
*+ bl_0_75 br_0_75 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c75
*+ bl_0_75 br_0_75 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c75
*+ bl_0_75 br_0_75 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c75
*+ bl_0_75 br_0_75 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c75
*+ bl_0_75 br_0_75 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c75
*+ bl_0_75 br_0_75 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c75
*+ bl_0_75 br_0_75 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c75
*+ bl_0_75 br_0_75 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c75
*+ bl_0_75 br_0_75 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c75
*+ bl_0_75 br_0_75 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c75
*+ bl_0_75 br_0_75 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c75
*+ bl_0_75 br_0_75 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c75
*+ bl_0_75 br_0_75 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c75
*+ bl_0_75 br_0_75 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c75
*+ bl_0_75 br_0_75 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c75
*+ bl_0_75 br_0_75 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c75
*+ bl_0_75 br_0_75 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c75
*+ bl_0_75 br_0_75 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c75
*+ bl_0_75 br_0_75 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c75
*+ bl_0_75 br_0_75 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c75
*+ bl_0_75 br_0_75 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c75
*+ bl_0_75 br_0_75 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c75
*+ bl_0_75 br_0_75 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c75
*+ bl_0_75 br_0_75 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c75
*+ bl_0_75 br_0_75 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c75
*+ bl_0_75 br_0_75 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c75
*+ bl_0_75 br_0_75 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c75
*+ bl_0_75 br_0_75 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c75
*+ bl_0_75 br_0_75 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c75
*+ bl_0_75 br_0_75 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c75
*+ bl_0_75 br_0_75 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c75
*+ bl_0_75 br_0_75 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c75
*+ bl_0_75 br_0_75 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c75
*+ bl_0_75 br_0_75 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c75
*+ bl_0_75 br_0_75 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c75
*+ bl_0_75 br_0_75 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c75
*+ bl_0_75 br_0_75 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c75
*+ bl_0_75 br_0_75 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c75
*+ bl_0_75 br_0_75 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c75
*+ bl_0_75 br_0_75 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c75
*+ bl_0_75 br_0_75 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c75
*+ bl_0_75 br_0_75 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c75
*+ bl_0_75 br_0_75 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c75
*+ bl_0_75 br_0_75 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c75
*+ bl_0_75 br_0_75 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c75
*+ bl_0_75 br_0_75 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c75
*+ bl_0_75 br_0_75 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c75
*+ bl_0_75 br_0_75 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c75
*+ bl_0_75 br_0_75 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c75
*+ bl_0_75 br_0_75 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c75
*+ bl_0_75 br_0_75 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c75
*+ bl_0_75 br_0_75 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c75
*+ bl_0_75 br_0_75 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c75
*+ bl_0_75 br_0_75 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c75
*+ bl_0_75 br_0_75 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c75
*+ bl_0_75 br_0_75 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c75
*+ bl_0_75 br_0_75 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c75
*+ bl_0_75 br_0_75 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c75
*+ bl_0_75 br_0_75 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c75
*+ bl_0_75 br_0_75 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c75
*+ bl_0_75 br_0_75 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c75
*+ bl_0_75 br_0_75 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c75
*+ bl_0_75 br_0_75 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c75
*+ bl_0_75 br_0_75 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c75
*+ bl_0_75 br_0_75 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c75
*+ bl_0_75 br_0_75 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c75
*+ bl_0_75 br_0_75 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c75
*+ bl_0_75 br_0_75 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c75
*+ bl_0_75 br_0_75 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c75
*+ bl_0_75 br_0_75 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c75
*+ bl_0_75 br_0_75 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c75
*+ bl_0_75 br_0_75 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c75
*+ bl_0_75 br_0_75 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c75
*+ bl_0_75 br_0_75 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c75
*+ bl_0_75 br_0_75 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c75
*+ bl_0_75 br_0_75 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c75
*+ bl_0_75 br_0_75 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c75
*+ bl_0_75 br_0_75 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c75
*+ bl_0_75 br_0_75 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c75
*+ bl_0_75 br_0_75 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c75
*+ bl_0_75 br_0_75 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c75
*+ bl_0_75 br_0_75 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c75
*+ bl_0_75 br_0_75 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c75
*+ bl_0_75 br_0_75 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c75
*+ bl_0_75 br_0_75 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c75
*+ bl_0_75 br_0_75 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c75
*+ bl_0_75 br_0_75 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c75
*+ bl_0_75 br_0_75 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c75
*+ bl_0_75 br_0_75 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c75
*+ bl_0_75 br_0_75 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c75
*+ bl_0_75 br_0_75 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c75
+ bl_0_75 br_0_75 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c76
+ bl_0_76 br_0_76 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c76
*+ bl_0_76 br_0_76 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c76
*+ bl_0_76 br_0_76 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c76
*+ bl_0_76 br_0_76 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c76
*+ bl_0_76 br_0_76 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c76
*+ bl_0_76 br_0_76 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c76
*+ bl_0_76 br_0_76 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c76
*+ bl_0_76 br_0_76 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c76
*+ bl_0_76 br_0_76 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c76
*+ bl_0_76 br_0_76 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c76
*+ bl_0_76 br_0_76 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c76
*+ bl_0_76 br_0_76 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c76
*+ bl_0_76 br_0_76 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c76
*+ bl_0_76 br_0_76 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c76
*+ bl_0_76 br_0_76 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c76
*+ bl_0_76 br_0_76 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c76
*+ bl_0_76 br_0_76 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c76
*+ bl_0_76 br_0_76 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c76
*+ bl_0_76 br_0_76 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c76
*+ bl_0_76 br_0_76 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c76
*+ bl_0_76 br_0_76 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c76
*+ bl_0_76 br_0_76 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c76
*+ bl_0_76 br_0_76 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c76
*+ bl_0_76 br_0_76 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c76
*+ bl_0_76 br_0_76 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c76
*+ bl_0_76 br_0_76 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c76
*+ bl_0_76 br_0_76 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c76
*+ bl_0_76 br_0_76 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c76
*+ bl_0_76 br_0_76 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c76
*+ bl_0_76 br_0_76 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c76
*+ bl_0_76 br_0_76 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c76
*+ bl_0_76 br_0_76 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c76
*+ bl_0_76 br_0_76 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c76
*+ bl_0_76 br_0_76 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c76
*+ bl_0_76 br_0_76 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c76
*+ bl_0_76 br_0_76 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c76
*+ bl_0_76 br_0_76 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c76
*+ bl_0_76 br_0_76 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c76
*+ bl_0_76 br_0_76 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c76
*+ bl_0_76 br_0_76 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c76
*+ bl_0_76 br_0_76 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c76
*+ bl_0_76 br_0_76 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c76
*+ bl_0_76 br_0_76 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c76
*+ bl_0_76 br_0_76 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c76
*+ bl_0_76 br_0_76 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c76
*+ bl_0_76 br_0_76 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c76
*+ bl_0_76 br_0_76 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c76
*+ bl_0_76 br_0_76 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c76
*+ bl_0_76 br_0_76 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c76
*+ bl_0_76 br_0_76 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c76
*+ bl_0_76 br_0_76 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c76
*+ bl_0_76 br_0_76 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c76
*+ bl_0_76 br_0_76 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c76
*+ bl_0_76 br_0_76 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c76
*+ bl_0_76 br_0_76 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c76
*+ bl_0_76 br_0_76 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c76
*+ bl_0_76 br_0_76 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c76
*+ bl_0_76 br_0_76 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c76
*+ bl_0_76 br_0_76 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c76
*+ bl_0_76 br_0_76 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c76
*+ bl_0_76 br_0_76 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c76
*+ bl_0_76 br_0_76 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c76
*+ bl_0_76 br_0_76 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c76
*+ bl_0_76 br_0_76 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c76
*+ bl_0_76 br_0_76 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c76
*+ bl_0_76 br_0_76 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c76
*+ bl_0_76 br_0_76 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c76
*+ bl_0_76 br_0_76 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c76
*+ bl_0_76 br_0_76 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c76
*+ bl_0_76 br_0_76 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c76
*+ bl_0_76 br_0_76 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c76
*+ bl_0_76 br_0_76 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c76
*+ bl_0_76 br_0_76 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c76
*+ bl_0_76 br_0_76 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c76
*+ bl_0_76 br_0_76 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c76
*+ bl_0_76 br_0_76 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c76
*+ bl_0_76 br_0_76 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c76
*+ bl_0_76 br_0_76 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c76
*+ bl_0_76 br_0_76 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c76
*+ bl_0_76 br_0_76 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c76
*+ bl_0_76 br_0_76 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c76
*+ bl_0_76 br_0_76 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c76
*+ bl_0_76 br_0_76 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c76
*+ bl_0_76 br_0_76 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c76
*+ bl_0_76 br_0_76 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c76
*+ bl_0_76 br_0_76 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c76
*+ bl_0_76 br_0_76 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c76
*+ bl_0_76 br_0_76 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c76
*+ bl_0_76 br_0_76 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c76
*+ bl_0_76 br_0_76 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c76
*+ bl_0_76 br_0_76 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c76
*+ bl_0_76 br_0_76 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c76
*+ bl_0_76 br_0_76 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c76
*+ bl_0_76 br_0_76 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c76
*+ bl_0_76 br_0_76 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c76
*+ bl_0_76 br_0_76 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c76
*+ bl_0_76 br_0_76 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c76
*+ bl_0_76 br_0_76 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c76
*+ bl_0_76 br_0_76 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c76
*+ bl_0_76 br_0_76 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c76
*+ bl_0_76 br_0_76 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c76
*+ bl_0_76 br_0_76 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c76
*+ bl_0_76 br_0_76 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c76
*+ bl_0_76 br_0_76 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c76
*+ bl_0_76 br_0_76 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c76
*+ bl_0_76 br_0_76 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c76
*+ bl_0_76 br_0_76 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c76
*+ bl_0_76 br_0_76 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c76
*+ bl_0_76 br_0_76 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c76
*+ bl_0_76 br_0_76 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c76
*+ bl_0_76 br_0_76 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c76
*+ bl_0_76 br_0_76 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c76
*+ bl_0_76 br_0_76 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c76
*+ bl_0_76 br_0_76 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c76
*+ bl_0_76 br_0_76 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c76
*+ bl_0_76 br_0_76 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c76
*+ bl_0_76 br_0_76 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c76
*+ bl_0_76 br_0_76 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c76
*+ bl_0_76 br_0_76 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c76
*+ bl_0_76 br_0_76 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c76
*+ bl_0_76 br_0_76 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c76
*+ bl_0_76 br_0_76 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c76
*+ bl_0_76 br_0_76 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c76
*+ bl_0_76 br_0_76 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c76
*+ bl_0_76 br_0_76 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c76
*+ bl_0_76 br_0_76 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c76
*+ bl_0_76 br_0_76 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c76
+ bl_0_76 br_0_76 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c77
+ bl_0_77 br_0_77 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c77
*+ bl_0_77 br_0_77 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c77
*+ bl_0_77 br_0_77 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c77
*+ bl_0_77 br_0_77 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c77
*+ bl_0_77 br_0_77 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c77
*+ bl_0_77 br_0_77 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c77
*+ bl_0_77 br_0_77 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c77
*+ bl_0_77 br_0_77 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c77
*+ bl_0_77 br_0_77 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c77
*+ bl_0_77 br_0_77 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c77
*+ bl_0_77 br_0_77 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c77
*+ bl_0_77 br_0_77 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c77
*+ bl_0_77 br_0_77 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c77
*+ bl_0_77 br_0_77 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c77
*+ bl_0_77 br_0_77 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c77
*+ bl_0_77 br_0_77 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c77
*+ bl_0_77 br_0_77 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c77
*+ bl_0_77 br_0_77 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c77
*+ bl_0_77 br_0_77 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c77
*+ bl_0_77 br_0_77 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c77
*+ bl_0_77 br_0_77 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c77
*+ bl_0_77 br_0_77 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c77
*+ bl_0_77 br_0_77 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c77
*+ bl_0_77 br_0_77 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c77
*+ bl_0_77 br_0_77 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c77
*+ bl_0_77 br_0_77 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c77
*+ bl_0_77 br_0_77 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c77
*+ bl_0_77 br_0_77 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c77
*+ bl_0_77 br_0_77 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c77
*+ bl_0_77 br_0_77 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c77
*+ bl_0_77 br_0_77 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c77
*+ bl_0_77 br_0_77 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c77
*+ bl_0_77 br_0_77 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c77
*+ bl_0_77 br_0_77 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c77
*+ bl_0_77 br_0_77 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c77
*+ bl_0_77 br_0_77 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c77
*+ bl_0_77 br_0_77 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c77
*+ bl_0_77 br_0_77 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c77
*+ bl_0_77 br_0_77 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c77
*+ bl_0_77 br_0_77 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c77
*+ bl_0_77 br_0_77 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c77
*+ bl_0_77 br_0_77 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c77
*+ bl_0_77 br_0_77 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c77
*+ bl_0_77 br_0_77 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c77
*+ bl_0_77 br_0_77 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c77
*+ bl_0_77 br_0_77 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c77
*+ bl_0_77 br_0_77 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c77
*+ bl_0_77 br_0_77 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c77
*+ bl_0_77 br_0_77 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c77
*+ bl_0_77 br_0_77 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c77
*+ bl_0_77 br_0_77 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c77
*+ bl_0_77 br_0_77 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c77
*+ bl_0_77 br_0_77 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c77
*+ bl_0_77 br_0_77 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c77
*+ bl_0_77 br_0_77 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c77
*+ bl_0_77 br_0_77 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c77
*+ bl_0_77 br_0_77 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c77
*+ bl_0_77 br_0_77 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c77
*+ bl_0_77 br_0_77 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c77
*+ bl_0_77 br_0_77 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c77
*+ bl_0_77 br_0_77 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c77
*+ bl_0_77 br_0_77 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c77
*+ bl_0_77 br_0_77 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c77
*+ bl_0_77 br_0_77 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c77
*+ bl_0_77 br_0_77 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c77
*+ bl_0_77 br_0_77 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c77
*+ bl_0_77 br_0_77 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c77
*+ bl_0_77 br_0_77 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c77
*+ bl_0_77 br_0_77 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c77
*+ bl_0_77 br_0_77 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c77
*+ bl_0_77 br_0_77 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c77
*+ bl_0_77 br_0_77 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c77
*+ bl_0_77 br_0_77 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c77
*+ bl_0_77 br_0_77 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c77
*+ bl_0_77 br_0_77 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c77
*+ bl_0_77 br_0_77 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c77
*+ bl_0_77 br_0_77 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c77
*+ bl_0_77 br_0_77 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c77
*+ bl_0_77 br_0_77 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c77
*+ bl_0_77 br_0_77 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c77
*+ bl_0_77 br_0_77 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c77
*+ bl_0_77 br_0_77 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c77
*+ bl_0_77 br_0_77 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c77
*+ bl_0_77 br_0_77 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c77
*+ bl_0_77 br_0_77 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c77
*+ bl_0_77 br_0_77 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c77
*+ bl_0_77 br_0_77 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c77
*+ bl_0_77 br_0_77 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c77
*+ bl_0_77 br_0_77 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c77
*+ bl_0_77 br_0_77 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c77
*+ bl_0_77 br_0_77 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c77
*+ bl_0_77 br_0_77 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c77
*+ bl_0_77 br_0_77 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c77
*+ bl_0_77 br_0_77 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c77
*+ bl_0_77 br_0_77 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c77
*+ bl_0_77 br_0_77 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c77
*+ bl_0_77 br_0_77 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c77
*+ bl_0_77 br_0_77 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c77
*+ bl_0_77 br_0_77 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c77
*+ bl_0_77 br_0_77 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c77
*+ bl_0_77 br_0_77 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c77
*+ bl_0_77 br_0_77 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c77
*+ bl_0_77 br_0_77 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c77
*+ bl_0_77 br_0_77 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c77
*+ bl_0_77 br_0_77 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c77
*+ bl_0_77 br_0_77 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c77
*+ bl_0_77 br_0_77 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c77
*+ bl_0_77 br_0_77 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c77
*+ bl_0_77 br_0_77 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c77
*+ bl_0_77 br_0_77 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c77
*+ bl_0_77 br_0_77 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c77
*+ bl_0_77 br_0_77 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c77
*+ bl_0_77 br_0_77 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c77
*+ bl_0_77 br_0_77 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c77
*+ bl_0_77 br_0_77 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c77
*+ bl_0_77 br_0_77 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c77
*+ bl_0_77 br_0_77 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c77
*+ bl_0_77 br_0_77 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c77
*+ bl_0_77 br_0_77 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c77
*+ bl_0_77 br_0_77 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c77
*+ bl_0_77 br_0_77 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c77
*+ bl_0_77 br_0_77 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c77
*+ bl_0_77 br_0_77 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c77
*+ bl_0_77 br_0_77 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c77
*+ bl_0_77 br_0_77 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c77
*+ bl_0_77 br_0_77 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c77
*+ bl_0_77 br_0_77 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c77
+ bl_0_77 br_0_77 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c78
+ bl_0_78 br_0_78 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c78
*+ bl_0_78 br_0_78 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c78
*+ bl_0_78 br_0_78 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c78
*+ bl_0_78 br_0_78 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c78
*+ bl_0_78 br_0_78 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c78
*+ bl_0_78 br_0_78 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c78
*+ bl_0_78 br_0_78 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c78
*+ bl_0_78 br_0_78 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c78
*+ bl_0_78 br_0_78 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c78
*+ bl_0_78 br_0_78 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c78
*+ bl_0_78 br_0_78 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c78
*+ bl_0_78 br_0_78 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c78
*+ bl_0_78 br_0_78 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c78
*+ bl_0_78 br_0_78 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c78
*+ bl_0_78 br_0_78 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c78
*+ bl_0_78 br_0_78 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c78
*+ bl_0_78 br_0_78 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c78
*+ bl_0_78 br_0_78 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c78
*+ bl_0_78 br_0_78 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c78
*+ bl_0_78 br_0_78 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c78
*+ bl_0_78 br_0_78 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c78
*+ bl_0_78 br_0_78 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c78
*+ bl_0_78 br_0_78 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c78
*+ bl_0_78 br_0_78 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c78
*+ bl_0_78 br_0_78 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c78
*+ bl_0_78 br_0_78 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c78
*+ bl_0_78 br_0_78 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c78
*+ bl_0_78 br_0_78 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c78
*+ bl_0_78 br_0_78 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c78
*+ bl_0_78 br_0_78 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c78
*+ bl_0_78 br_0_78 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c78
*+ bl_0_78 br_0_78 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c78
*+ bl_0_78 br_0_78 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c78
*+ bl_0_78 br_0_78 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c78
*+ bl_0_78 br_0_78 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c78
*+ bl_0_78 br_0_78 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c78
*+ bl_0_78 br_0_78 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c78
*+ bl_0_78 br_0_78 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c78
*+ bl_0_78 br_0_78 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c78
*+ bl_0_78 br_0_78 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c78
*+ bl_0_78 br_0_78 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c78
*+ bl_0_78 br_0_78 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c78
*+ bl_0_78 br_0_78 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c78
*+ bl_0_78 br_0_78 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c78
*+ bl_0_78 br_0_78 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c78
*+ bl_0_78 br_0_78 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c78
*+ bl_0_78 br_0_78 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c78
*+ bl_0_78 br_0_78 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c78
*+ bl_0_78 br_0_78 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c78
*+ bl_0_78 br_0_78 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c78
*+ bl_0_78 br_0_78 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c78
*+ bl_0_78 br_0_78 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c78
*+ bl_0_78 br_0_78 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c78
*+ bl_0_78 br_0_78 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c78
*+ bl_0_78 br_0_78 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c78
*+ bl_0_78 br_0_78 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c78
*+ bl_0_78 br_0_78 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c78
*+ bl_0_78 br_0_78 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c78
*+ bl_0_78 br_0_78 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c78
*+ bl_0_78 br_0_78 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c78
*+ bl_0_78 br_0_78 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c78
*+ bl_0_78 br_0_78 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c78
*+ bl_0_78 br_0_78 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c78
*+ bl_0_78 br_0_78 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c78
*+ bl_0_78 br_0_78 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c78
*+ bl_0_78 br_0_78 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c78
*+ bl_0_78 br_0_78 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c78
*+ bl_0_78 br_0_78 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c78
*+ bl_0_78 br_0_78 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c78
*+ bl_0_78 br_0_78 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c78
*+ bl_0_78 br_0_78 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c78
*+ bl_0_78 br_0_78 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c78
*+ bl_0_78 br_0_78 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c78
*+ bl_0_78 br_0_78 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c78
*+ bl_0_78 br_0_78 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c78
*+ bl_0_78 br_0_78 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c78
*+ bl_0_78 br_0_78 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c78
*+ bl_0_78 br_0_78 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c78
*+ bl_0_78 br_0_78 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c78
*+ bl_0_78 br_0_78 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c78
*+ bl_0_78 br_0_78 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c78
*+ bl_0_78 br_0_78 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c78
*+ bl_0_78 br_0_78 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c78
*+ bl_0_78 br_0_78 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c78
*+ bl_0_78 br_0_78 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c78
*+ bl_0_78 br_0_78 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c78
*+ bl_0_78 br_0_78 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c78
*+ bl_0_78 br_0_78 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c78
*+ bl_0_78 br_0_78 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c78
*+ bl_0_78 br_0_78 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c78
*+ bl_0_78 br_0_78 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c78
*+ bl_0_78 br_0_78 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c78
*+ bl_0_78 br_0_78 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c78
*+ bl_0_78 br_0_78 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c78
*+ bl_0_78 br_0_78 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c78
*+ bl_0_78 br_0_78 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c78
*+ bl_0_78 br_0_78 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c78
*+ bl_0_78 br_0_78 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c78
*+ bl_0_78 br_0_78 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c78
*+ bl_0_78 br_0_78 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c78
*+ bl_0_78 br_0_78 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c78
*+ bl_0_78 br_0_78 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c78
*+ bl_0_78 br_0_78 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c78
*+ bl_0_78 br_0_78 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c78
*+ bl_0_78 br_0_78 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c78
*+ bl_0_78 br_0_78 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c78
*+ bl_0_78 br_0_78 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c78
*+ bl_0_78 br_0_78 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c78
*+ bl_0_78 br_0_78 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c78
*+ bl_0_78 br_0_78 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c78
*+ bl_0_78 br_0_78 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c78
*+ bl_0_78 br_0_78 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c78
*+ bl_0_78 br_0_78 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c78
*+ bl_0_78 br_0_78 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c78
*+ bl_0_78 br_0_78 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c78
*+ bl_0_78 br_0_78 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c78
*+ bl_0_78 br_0_78 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c78
*+ bl_0_78 br_0_78 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c78
*+ bl_0_78 br_0_78 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c78
*+ bl_0_78 br_0_78 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c78
*+ bl_0_78 br_0_78 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c78
*+ bl_0_78 br_0_78 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c78
*+ bl_0_78 br_0_78 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c78
*+ bl_0_78 br_0_78 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c78
*+ bl_0_78 br_0_78 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c78
*+ bl_0_78 br_0_78 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c78
*+ bl_0_78 br_0_78 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c78
+ bl_0_78 br_0_78 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c79
+ bl_0_79 br_0_79 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c79
*+ bl_0_79 br_0_79 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c79
*+ bl_0_79 br_0_79 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c79
*+ bl_0_79 br_0_79 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c79
*+ bl_0_79 br_0_79 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c79
*+ bl_0_79 br_0_79 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c79
*+ bl_0_79 br_0_79 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c79
*+ bl_0_79 br_0_79 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c79
*+ bl_0_79 br_0_79 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c79
*+ bl_0_79 br_0_79 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c79
*+ bl_0_79 br_0_79 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c79
*+ bl_0_79 br_0_79 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c79
*+ bl_0_79 br_0_79 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c79
*+ bl_0_79 br_0_79 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c79
*+ bl_0_79 br_0_79 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c79
*+ bl_0_79 br_0_79 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c79
*+ bl_0_79 br_0_79 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c79
*+ bl_0_79 br_0_79 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c79
*+ bl_0_79 br_0_79 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c79
*+ bl_0_79 br_0_79 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c79
*+ bl_0_79 br_0_79 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c79
*+ bl_0_79 br_0_79 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c79
*+ bl_0_79 br_0_79 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c79
*+ bl_0_79 br_0_79 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c79
*+ bl_0_79 br_0_79 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c79
*+ bl_0_79 br_0_79 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c79
*+ bl_0_79 br_0_79 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c79
*+ bl_0_79 br_0_79 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c79
*+ bl_0_79 br_0_79 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c79
*+ bl_0_79 br_0_79 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c79
*+ bl_0_79 br_0_79 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c79
*+ bl_0_79 br_0_79 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c79
*+ bl_0_79 br_0_79 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c79
*+ bl_0_79 br_0_79 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c79
*+ bl_0_79 br_0_79 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c79
*+ bl_0_79 br_0_79 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c79
*+ bl_0_79 br_0_79 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c79
*+ bl_0_79 br_0_79 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c79
*+ bl_0_79 br_0_79 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c79
*+ bl_0_79 br_0_79 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c79
*+ bl_0_79 br_0_79 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c79
*+ bl_0_79 br_0_79 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c79
*+ bl_0_79 br_0_79 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c79
*+ bl_0_79 br_0_79 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c79
*+ bl_0_79 br_0_79 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c79
*+ bl_0_79 br_0_79 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c79
*+ bl_0_79 br_0_79 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c79
*+ bl_0_79 br_0_79 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c79
*+ bl_0_79 br_0_79 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c79
*+ bl_0_79 br_0_79 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c79
*+ bl_0_79 br_0_79 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c79
*+ bl_0_79 br_0_79 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c79
*+ bl_0_79 br_0_79 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c79
*+ bl_0_79 br_0_79 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c79
*+ bl_0_79 br_0_79 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c79
*+ bl_0_79 br_0_79 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c79
*+ bl_0_79 br_0_79 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c79
*+ bl_0_79 br_0_79 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c79
*+ bl_0_79 br_0_79 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c79
*+ bl_0_79 br_0_79 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c79
*+ bl_0_79 br_0_79 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c79
*+ bl_0_79 br_0_79 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c79
*+ bl_0_79 br_0_79 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c79
*+ bl_0_79 br_0_79 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c79
*+ bl_0_79 br_0_79 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c79
*+ bl_0_79 br_0_79 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c79
*+ bl_0_79 br_0_79 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c79
*+ bl_0_79 br_0_79 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c79
*+ bl_0_79 br_0_79 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c79
*+ bl_0_79 br_0_79 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c79
*+ bl_0_79 br_0_79 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c79
*+ bl_0_79 br_0_79 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c79
*+ bl_0_79 br_0_79 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c79
*+ bl_0_79 br_0_79 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c79
*+ bl_0_79 br_0_79 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c79
*+ bl_0_79 br_0_79 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c79
*+ bl_0_79 br_0_79 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c79
*+ bl_0_79 br_0_79 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c79
*+ bl_0_79 br_0_79 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c79
*+ bl_0_79 br_0_79 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c79
*+ bl_0_79 br_0_79 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c79
*+ bl_0_79 br_0_79 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c79
*+ bl_0_79 br_0_79 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c79
*+ bl_0_79 br_0_79 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c79
*+ bl_0_79 br_0_79 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c79
*+ bl_0_79 br_0_79 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c79
*+ bl_0_79 br_0_79 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c79
*+ bl_0_79 br_0_79 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c79
*+ bl_0_79 br_0_79 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c79
*+ bl_0_79 br_0_79 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c79
*+ bl_0_79 br_0_79 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c79
*+ bl_0_79 br_0_79 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c79
*+ bl_0_79 br_0_79 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c79
*+ bl_0_79 br_0_79 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c79
*+ bl_0_79 br_0_79 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c79
*+ bl_0_79 br_0_79 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c79
*+ bl_0_79 br_0_79 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c79
*+ bl_0_79 br_0_79 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c79
*+ bl_0_79 br_0_79 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c79
*+ bl_0_79 br_0_79 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c79
*+ bl_0_79 br_0_79 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c79
*+ bl_0_79 br_0_79 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c79
*+ bl_0_79 br_0_79 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c79
*+ bl_0_79 br_0_79 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c79
*+ bl_0_79 br_0_79 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c79
*+ bl_0_79 br_0_79 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c79
*+ bl_0_79 br_0_79 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c79
*+ bl_0_79 br_0_79 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c79
*+ bl_0_79 br_0_79 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c79
*+ bl_0_79 br_0_79 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c79
*+ bl_0_79 br_0_79 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c79
*+ bl_0_79 br_0_79 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c79
*+ bl_0_79 br_0_79 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c79
*+ bl_0_79 br_0_79 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c79
*+ bl_0_79 br_0_79 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c79
*+ bl_0_79 br_0_79 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c79
*+ bl_0_79 br_0_79 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c79
*+ bl_0_79 br_0_79 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c79
*+ bl_0_79 br_0_79 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c79
*+ bl_0_79 br_0_79 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c79
*+ bl_0_79 br_0_79 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c79
*+ bl_0_79 br_0_79 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c79
*+ bl_0_79 br_0_79 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c79
*+ bl_0_79 br_0_79 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c79
*+ bl_0_79 br_0_79 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c79
*+ bl_0_79 br_0_79 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c79
*+ bl_0_79 br_0_79 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c79
+ bl_0_79 br_0_79 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c80
+ bl_0_80 br_0_80 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c80
*+ bl_0_80 br_0_80 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c80
*+ bl_0_80 br_0_80 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c80
*+ bl_0_80 br_0_80 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c80
*+ bl_0_80 br_0_80 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c80
*+ bl_0_80 br_0_80 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c80
*+ bl_0_80 br_0_80 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c80
*+ bl_0_80 br_0_80 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c80
*+ bl_0_80 br_0_80 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c80
*+ bl_0_80 br_0_80 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c80
*+ bl_0_80 br_0_80 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c80
*+ bl_0_80 br_0_80 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c80
*+ bl_0_80 br_0_80 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c80
*+ bl_0_80 br_0_80 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c80
*+ bl_0_80 br_0_80 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c80
*+ bl_0_80 br_0_80 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c80
*+ bl_0_80 br_0_80 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c80
*+ bl_0_80 br_0_80 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c80
*+ bl_0_80 br_0_80 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c80
*+ bl_0_80 br_0_80 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c80
*+ bl_0_80 br_0_80 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c80
*+ bl_0_80 br_0_80 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c80
*+ bl_0_80 br_0_80 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c80
*+ bl_0_80 br_0_80 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c80
*+ bl_0_80 br_0_80 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c80
*+ bl_0_80 br_0_80 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c80
*+ bl_0_80 br_0_80 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c80
*+ bl_0_80 br_0_80 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c80
*+ bl_0_80 br_0_80 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c80
*+ bl_0_80 br_0_80 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c80
*+ bl_0_80 br_0_80 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c80
*+ bl_0_80 br_0_80 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c80
*+ bl_0_80 br_0_80 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c80
*+ bl_0_80 br_0_80 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c80
*+ bl_0_80 br_0_80 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c80
*+ bl_0_80 br_0_80 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c80
*+ bl_0_80 br_0_80 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c80
*+ bl_0_80 br_0_80 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c80
*+ bl_0_80 br_0_80 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c80
*+ bl_0_80 br_0_80 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c80
*+ bl_0_80 br_0_80 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c80
*+ bl_0_80 br_0_80 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c80
*+ bl_0_80 br_0_80 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c80
*+ bl_0_80 br_0_80 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c80
*+ bl_0_80 br_0_80 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c80
*+ bl_0_80 br_0_80 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c80
*+ bl_0_80 br_0_80 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c80
*+ bl_0_80 br_0_80 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c80
*+ bl_0_80 br_0_80 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c80
*+ bl_0_80 br_0_80 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c80
*+ bl_0_80 br_0_80 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c80
*+ bl_0_80 br_0_80 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c80
*+ bl_0_80 br_0_80 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c80
*+ bl_0_80 br_0_80 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c80
*+ bl_0_80 br_0_80 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c80
*+ bl_0_80 br_0_80 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c80
*+ bl_0_80 br_0_80 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c80
*+ bl_0_80 br_0_80 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c80
*+ bl_0_80 br_0_80 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c80
*+ bl_0_80 br_0_80 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c80
*+ bl_0_80 br_0_80 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c80
*+ bl_0_80 br_0_80 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c80
*+ bl_0_80 br_0_80 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c80
*+ bl_0_80 br_0_80 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c80
*+ bl_0_80 br_0_80 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c80
*+ bl_0_80 br_0_80 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c80
*+ bl_0_80 br_0_80 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c80
*+ bl_0_80 br_0_80 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c80
*+ bl_0_80 br_0_80 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c80
*+ bl_0_80 br_0_80 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c80
*+ bl_0_80 br_0_80 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c80
*+ bl_0_80 br_0_80 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c80
*+ bl_0_80 br_0_80 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c80
*+ bl_0_80 br_0_80 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c80
*+ bl_0_80 br_0_80 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c80
*+ bl_0_80 br_0_80 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c80
*+ bl_0_80 br_0_80 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c80
*+ bl_0_80 br_0_80 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c80
*+ bl_0_80 br_0_80 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c80
*+ bl_0_80 br_0_80 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c80
*+ bl_0_80 br_0_80 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c80
*+ bl_0_80 br_0_80 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c80
*+ bl_0_80 br_0_80 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c80
*+ bl_0_80 br_0_80 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c80
*+ bl_0_80 br_0_80 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c80
*+ bl_0_80 br_0_80 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c80
*+ bl_0_80 br_0_80 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c80
*+ bl_0_80 br_0_80 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c80
*+ bl_0_80 br_0_80 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c80
*+ bl_0_80 br_0_80 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c80
*+ bl_0_80 br_0_80 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c80
*+ bl_0_80 br_0_80 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c80
*+ bl_0_80 br_0_80 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c80
*+ bl_0_80 br_0_80 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c80
*+ bl_0_80 br_0_80 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c80
*+ bl_0_80 br_0_80 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c80
*+ bl_0_80 br_0_80 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c80
*+ bl_0_80 br_0_80 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c80
*+ bl_0_80 br_0_80 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c80
*+ bl_0_80 br_0_80 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c80
*+ bl_0_80 br_0_80 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c80
*+ bl_0_80 br_0_80 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c80
*+ bl_0_80 br_0_80 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c80
*+ bl_0_80 br_0_80 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c80
*+ bl_0_80 br_0_80 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c80
*+ bl_0_80 br_0_80 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c80
*+ bl_0_80 br_0_80 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c80
*+ bl_0_80 br_0_80 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c80
*+ bl_0_80 br_0_80 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c80
*+ bl_0_80 br_0_80 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c80
*+ bl_0_80 br_0_80 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c80
*+ bl_0_80 br_0_80 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c80
*+ bl_0_80 br_0_80 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c80
*+ bl_0_80 br_0_80 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c80
*+ bl_0_80 br_0_80 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c80
*+ bl_0_80 br_0_80 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c80
*+ bl_0_80 br_0_80 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c80
*+ bl_0_80 br_0_80 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c80
*+ bl_0_80 br_0_80 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c80
*+ bl_0_80 br_0_80 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c80
*+ bl_0_80 br_0_80 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c80
*+ bl_0_80 br_0_80 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c80
*+ bl_0_80 br_0_80 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c80
*+ bl_0_80 br_0_80 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c80
*+ bl_0_80 br_0_80 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c80
*+ bl_0_80 br_0_80 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c80
*+ bl_0_80 br_0_80 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c80
+ bl_0_80 br_0_80 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c81
+ bl_0_81 br_0_81 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c81
*+ bl_0_81 br_0_81 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c81
*+ bl_0_81 br_0_81 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c81
*+ bl_0_81 br_0_81 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c81
*+ bl_0_81 br_0_81 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c81
*+ bl_0_81 br_0_81 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c81
*+ bl_0_81 br_0_81 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c81
*+ bl_0_81 br_0_81 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c81
*+ bl_0_81 br_0_81 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c81
*+ bl_0_81 br_0_81 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c81
*+ bl_0_81 br_0_81 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c81
*+ bl_0_81 br_0_81 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c81
*+ bl_0_81 br_0_81 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c81
*+ bl_0_81 br_0_81 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c81
*+ bl_0_81 br_0_81 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c81
*+ bl_0_81 br_0_81 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c81
*+ bl_0_81 br_0_81 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c81
*+ bl_0_81 br_0_81 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c81
*+ bl_0_81 br_0_81 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c81
*+ bl_0_81 br_0_81 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c81
*+ bl_0_81 br_0_81 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c81
*+ bl_0_81 br_0_81 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c81
*+ bl_0_81 br_0_81 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c81
*+ bl_0_81 br_0_81 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c81
*+ bl_0_81 br_0_81 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c81
*+ bl_0_81 br_0_81 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c81
*+ bl_0_81 br_0_81 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c81
*+ bl_0_81 br_0_81 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c81
*+ bl_0_81 br_0_81 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c81
*+ bl_0_81 br_0_81 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c81
*+ bl_0_81 br_0_81 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c81
*+ bl_0_81 br_0_81 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c81
*+ bl_0_81 br_0_81 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c81
*+ bl_0_81 br_0_81 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c81
*+ bl_0_81 br_0_81 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c81
*+ bl_0_81 br_0_81 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c81
*+ bl_0_81 br_0_81 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c81
*+ bl_0_81 br_0_81 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c81
*+ bl_0_81 br_0_81 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c81
*+ bl_0_81 br_0_81 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c81
*+ bl_0_81 br_0_81 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c81
*+ bl_0_81 br_0_81 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c81
*+ bl_0_81 br_0_81 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c81
*+ bl_0_81 br_0_81 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c81
*+ bl_0_81 br_0_81 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c81
*+ bl_0_81 br_0_81 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c81
*+ bl_0_81 br_0_81 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c81
*+ bl_0_81 br_0_81 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c81
*+ bl_0_81 br_0_81 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c81
*+ bl_0_81 br_0_81 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c81
*+ bl_0_81 br_0_81 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c81
*+ bl_0_81 br_0_81 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c81
*+ bl_0_81 br_0_81 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c81
*+ bl_0_81 br_0_81 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c81
*+ bl_0_81 br_0_81 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c81
*+ bl_0_81 br_0_81 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c81
*+ bl_0_81 br_0_81 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c81
*+ bl_0_81 br_0_81 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c81
*+ bl_0_81 br_0_81 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c81
*+ bl_0_81 br_0_81 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c81
*+ bl_0_81 br_0_81 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c81
*+ bl_0_81 br_0_81 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c81
*+ bl_0_81 br_0_81 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c81
*+ bl_0_81 br_0_81 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c81
*+ bl_0_81 br_0_81 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c81
*+ bl_0_81 br_0_81 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c81
*+ bl_0_81 br_0_81 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c81
*+ bl_0_81 br_0_81 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c81
*+ bl_0_81 br_0_81 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c81
*+ bl_0_81 br_0_81 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c81
*+ bl_0_81 br_0_81 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c81
*+ bl_0_81 br_0_81 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c81
*+ bl_0_81 br_0_81 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c81
*+ bl_0_81 br_0_81 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c81
*+ bl_0_81 br_0_81 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c81
*+ bl_0_81 br_0_81 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c81
*+ bl_0_81 br_0_81 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c81
*+ bl_0_81 br_0_81 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c81
*+ bl_0_81 br_0_81 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c81
*+ bl_0_81 br_0_81 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c81
*+ bl_0_81 br_0_81 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c81
*+ bl_0_81 br_0_81 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c81
*+ bl_0_81 br_0_81 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c81
*+ bl_0_81 br_0_81 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c81
*+ bl_0_81 br_0_81 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c81
*+ bl_0_81 br_0_81 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c81
*+ bl_0_81 br_0_81 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c81
*+ bl_0_81 br_0_81 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c81
*+ bl_0_81 br_0_81 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c81
*+ bl_0_81 br_0_81 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c81
*+ bl_0_81 br_0_81 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c81
*+ bl_0_81 br_0_81 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c81
*+ bl_0_81 br_0_81 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c81
*+ bl_0_81 br_0_81 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c81
*+ bl_0_81 br_0_81 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c81
*+ bl_0_81 br_0_81 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c81
*+ bl_0_81 br_0_81 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c81
*+ bl_0_81 br_0_81 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c81
*+ bl_0_81 br_0_81 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c81
*+ bl_0_81 br_0_81 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c81
*+ bl_0_81 br_0_81 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c81
*+ bl_0_81 br_0_81 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c81
*+ bl_0_81 br_0_81 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c81
*+ bl_0_81 br_0_81 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c81
*+ bl_0_81 br_0_81 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c81
*+ bl_0_81 br_0_81 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c81
*+ bl_0_81 br_0_81 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c81
*+ bl_0_81 br_0_81 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c81
*+ bl_0_81 br_0_81 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c81
*+ bl_0_81 br_0_81 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c81
*+ bl_0_81 br_0_81 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c81
*+ bl_0_81 br_0_81 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c81
*+ bl_0_81 br_0_81 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c81
*+ bl_0_81 br_0_81 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c81
*+ bl_0_81 br_0_81 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c81
*+ bl_0_81 br_0_81 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c81
*+ bl_0_81 br_0_81 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c81
*+ bl_0_81 br_0_81 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c81
*+ bl_0_81 br_0_81 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c81
*+ bl_0_81 br_0_81 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c81
*+ bl_0_81 br_0_81 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c81
*+ bl_0_81 br_0_81 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c81
*+ bl_0_81 br_0_81 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c81
*+ bl_0_81 br_0_81 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c81
*+ bl_0_81 br_0_81 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c81
*+ bl_0_81 br_0_81 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c81
*+ bl_0_81 br_0_81 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c81
+ bl_0_81 br_0_81 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c82
+ bl_0_82 br_0_82 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c82
*+ bl_0_82 br_0_82 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c82
*+ bl_0_82 br_0_82 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c82
*+ bl_0_82 br_0_82 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c82
*+ bl_0_82 br_0_82 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c82
*+ bl_0_82 br_0_82 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c82
*+ bl_0_82 br_0_82 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c82
*+ bl_0_82 br_0_82 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c82
*+ bl_0_82 br_0_82 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c82
*+ bl_0_82 br_0_82 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c82
*+ bl_0_82 br_0_82 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c82
*+ bl_0_82 br_0_82 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c82
*+ bl_0_82 br_0_82 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c82
*+ bl_0_82 br_0_82 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c82
*+ bl_0_82 br_0_82 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c82
*+ bl_0_82 br_0_82 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c82
*+ bl_0_82 br_0_82 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c82
*+ bl_0_82 br_0_82 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c82
*+ bl_0_82 br_0_82 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c82
*+ bl_0_82 br_0_82 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c82
*+ bl_0_82 br_0_82 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c82
*+ bl_0_82 br_0_82 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c82
*+ bl_0_82 br_0_82 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c82
*+ bl_0_82 br_0_82 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c82
*+ bl_0_82 br_0_82 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c82
*+ bl_0_82 br_0_82 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c82
*+ bl_0_82 br_0_82 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c82
*+ bl_0_82 br_0_82 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c82
*+ bl_0_82 br_0_82 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c82
*+ bl_0_82 br_0_82 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c82
*+ bl_0_82 br_0_82 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c82
*+ bl_0_82 br_0_82 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c82
*+ bl_0_82 br_0_82 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c82
*+ bl_0_82 br_0_82 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c82
*+ bl_0_82 br_0_82 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c82
*+ bl_0_82 br_0_82 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c82
*+ bl_0_82 br_0_82 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c82
*+ bl_0_82 br_0_82 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c82
*+ bl_0_82 br_0_82 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c82
*+ bl_0_82 br_0_82 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c82
*+ bl_0_82 br_0_82 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c82
*+ bl_0_82 br_0_82 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c82
*+ bl_0_82 br_0_82 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c82
*+ bl_0_82 br_0_82 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c82
*+ bl_0_82 br_0_82 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c82
*+ bl_0_82 br_0_82 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c82
*+ bl_0_82 br_0_82 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c82
*+ bl_0_82 br_0_82 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c82
*+ bl_0_82 br_0_82 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c82
*+ bl_0_82 br_0_82 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c82
*+ bl_0_82 br_0_82 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c82
*+ bl_0_82 br_0_82 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c82
*+ bl_0_82 br_0_82 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c82
*+ bl_0_82 br_0_82 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c82
*+ bl_0_82 br_0_82 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c82
*+ bl_0_82 br_0_82 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c82
*+ bl_0_82 br_0_82 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c82
*+ bl_0_82 br_0_82 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c82
*+ bl_0_82 br_0_82 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c82
*+ bl_0_82 br_0_82 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c82
*+ bl_0_82 br_0_82 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c82
*+ bl_0_82 br_0_82 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c82
*+ bl_0_82 br_0_82 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c82
*+ bl_0_82 br_0_82 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c82
*+ bl_0_82 br_0_82 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c82
*+ bl_0_82 br_0_82 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c82
*+ bl_0_82 br_0_82 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c82
*+ bl_0_82 br_0_82 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c82
*+ bl_0_82 br_0_82 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c82
*+ bl_0_82 br_0_82 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c82
*+ bl_0_82 br_0_82 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c82
*+ bl_0_82 br_0_82 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c82
*+ bl_0_82 br_0_82 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c82
*+ bl_0_82 br_0_82 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c82
*+ bl_0_82 br_0_82 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c82
*+ bl_0_82 br_0_82 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c82
*+ bl_0_82 br_0_82 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c82
*+ bl_0_82 br_0_82 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c82
*+ bl_0_82 br_0_82 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c82
*+ bl_0_82 br_0_82 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c82
*+ bl_0_82 br_0_82 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c82
*+ bl_0_82 br_0_82 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c82
*+ bl_0_82 br_0_82 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c82
*+ bl_0_82 br_0_82 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c82
*+ bl_0_82 br_0_82 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c82
*+ bl_0_82 br_0_82 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c82
*+ bl_0_82 br_0_82 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c82
*+ bl_0_82 br_0_82 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c82
*+ bl_0_82 br_0_82 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c82
*+ bl_0_82 br_0_82 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c82
*+ bl_0_82 br_0_82 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c82
*+ bl_0_82 br_0_82 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c82
*+ bl_0_82 br_0_82 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c82
*+ bl_0_82 br_0_82 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c82
*+ bl_0_82 br_0_82 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c82
*+ bl_0_82 br_0_82 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c82
*+ bl_0_82 br_0_82 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c82
*+ bl_0_82 br_0_82 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c82
*+ bl_0_82 br_0_82 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c82
*+ bl_0_82 br_0_82 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c82
*+ bl_0_82 br_0_82 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c82
*+ bl_0_82 br_0_82 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c82
*+ bl_0_82 br_0_82 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c82
*+ bl_0_82 br_0_82 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c82
*+ bl_0_82 br_0_82 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c82
*+ bl_0_82 br_0_82 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c82
*+ bl_0_82 br_0_82 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c82
*+ bl_0_82 br_0_82 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c82
*+ bl_0_82 br_0_82 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c82
*+ bl_0_82 br_0_82 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c82
*+ bl_0_82 br_0_82 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c82
*+ bl_0_82 br_0_82 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c82
*+ bl_0_82 br_0_82 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c82
*+ bl_0_82 br_0_82 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c82
*+ bl_0_82 br_0_82 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c82
*+ bl_0_82 br_0_82 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c82
*+ bl_0_82 br_0_82 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c82
*+ bl_0_82 br_0_82 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c82
*+ bl_0_82 br_0_82 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c82
*+ bl_0_82 br_0_82 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c82
*+ bl_0_82 br_0_82 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c82
*+ bl_0_82 br_0_82 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c82
*+ bl_0_82 br_0_82 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c82
*+ bl_0_82 br_0_82 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c82
*+ bl_0_82 br_0_82 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c82
*+ bl_0_82 br_0_82 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c82
*+ bl_0_82 br_0_82 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c82
+ bl_0_82 br_0_82 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c83
+ bl_0_83 br_0_83 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c83
*+ bl_0_83 br_0_83 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c83
*+ bl_0_83 br_0_83 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c83
*+ bl_0_83 br_0_83 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c83
*+ bl_0_83 br_0_83 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c83
*+ bl_0_83 br_0_83 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c83
*+ bl_0_83 br_0_83 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c83
*+ bl_0_83 br_0_83 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c83
*+ bl_0_83 br_0_83 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c83
*+ bl_0_83 br_0_83 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c83
*+ bl_0_83 br_0_83 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c83
*+ bl_0_83 br_0_83 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c83
*+ bl_0_83 br_0_83 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c83
*+ bl_0_83 br_0_83 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c83
*+ bl_0_83 br_0_83 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c83
*+ bl_0_83 br_0_83 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c83
*+ bl_0_83 br_0_83 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c83
*+ bl_0_83 br_0_83 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c83
*+ bl_0_83 br_0_83 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c83
*+ bl_0_83 br_0_83 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c83
*+ bl_0_83 br_0_83 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c83
*+ bl_0_83 br_0_83 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c83
*+ bl_0_83 br_0_83 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c83
*+ bl_0_83 br_0_83 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c83
*+ bl_0_83 br_0_83 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c83
*+ bl_0_83 br_0_83 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c83
*+ bl_0_83 br_0_83 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c83
*+ bl_0_83 br_0_83 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c83
*+ bl_0_83 br_0_83 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c83
*+ bl_0_83 br_0_83 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c83
*+ bl_0_83 br_0_83 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c83
*+ bl_0_83 br_0_83 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c83
*+ bl_0_83 br_0_83 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c83
*+ bl_0_83 br_0_83 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c83
*+ bl_0_83 br_0_83 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c83
*+ bl_0_83 br_0_83 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c83
*+ bl_0_83 br_0_83 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c83
*+ bl_0_83 br_0_83 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c83
*+ bl_0_83 br_0_83 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c83
*+ bl_0_83 br_0_83 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c83
*+ bl_0_83 br_0_83 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c83
*+ bl_0_83 br_0_83 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c83
*+ bl_0_83 br_0_83 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c83
*+ bl_0_83 br_0_83 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c83
*+ bl_0_83 br_0_83 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c83
*+ bl_0_83 br_0_83 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c83
*+ bl_0_83 br_0_83 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c83
*+ bl_0_83 br_0_83 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c83
*+ bl_0_83 br_0_83 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c83
*+ bl_0_83 br_0_83 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c83
*+ bl_0_83 br_0_83 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c83
*+ bl_0_83 br_0_83 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c83
*+ bl_0_83 br_0_83 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c83
*+ bl_0_83 br_0_83 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c83
*+ bl_0_83 br_0_83 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c83
*+ bl_0_83 br_0_83 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c83
*+ bl_0_83 br_0_83 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c83
*+ bl_0_83 br_0_83 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c83
*+ bl_0_83 br_0_83 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c83
*+ bl_0_83 br_0_83 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c83
*+ bl_0_83 br_0_83 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c83
*+ bl_0_83 br_0_83 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c83
*+ bl_0_83 br_0_83 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c83
*+ bl_0_83 br_0_83 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c83
*+ bl_0_83 br_0_83 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c83
*+ bl_0_83 br_0_83 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c83
*+ bl_0_83 br_0_83 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c83
*+ bl_0_83 br_0_83 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c83
*+ bl_0_83 br_0_83 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c83
*+ bl_0_83 br_0_83 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c83
*+ bl_0_83 br_0_83 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c83
*+ bl_0_83 br_0_83 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c83
*+ bl_0_83 br_0_83 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c83
*+ bl_0_83 br_0_83 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c83
*+ bl_0_83 br_0_83 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c83
*+ bl_0_83 br_0_83 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c83
*+ bl_0_83 br_0_83 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c83
*+ bl_0_83 br_0_83 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c83
*+ bl_0_83 br_0_83 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c83
*+ bl_0_83 br_0_83 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c83
*+ bl_0_83 br_0_83 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c83
*+ bl_0_83 br_0_83 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c83
*+ bl_0_83 br_0_83 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c83
*+ bl_0_83 br_0_83 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c83
*+ bl_0_83 br_0_83 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c83
*+ bl_0_83 br_0_83 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c83
*+ bl_0_83 br_0_83 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c83
*+ bl_0_83 br_0_83 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c83
*+ bl_0_83 br_0_83 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c83
*+ bl_0_83 br_0_83 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c83
*+ bl_0_83 br_0_83 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c83
*+ bl_0_83 br_0_83 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c83
*+ bl_0_83 br_0_83 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c83
*+ bl_0_83 br_0_83 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c83
*+ bl_0_83 br_0_83 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c83
*+ bl_0_83 br_0_83 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c83
*+ bl_0_83 br_0_83 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c83
*+ bl_0_83 br_0_83 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c83
*+ bl_0_83 br_0_83 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c83
*+ bl_0_83 br_0_83 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c83
*+ bl_0_83 br_0_83 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c83
*+ bl_0_83 br_0_83 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c83
*+ bl_0_83 br_0_83 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c83
*+ bl_0_83 br_0_83 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c83
*+ bl_0_83 br_0_83 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c83
*+ bl_0_83 br_0_83 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c83
*+ bl_0_83 br_0_83 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c83
*+ bl_0_83 br_0_83 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c83
*+ bl_0_83 br_0_83 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c83
*+ bl_0_83 br_0_83 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c83
*+ bl_0_83 br_0_83 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c83
*+ bl_0_83 br_0_83 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c83
*+ bl_0_83 br_0_83 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c83
*+ bl_0_83 br_0_83 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c83
*+ bl_0_83 br_0_83 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c83
*+ bl_0_83 br_0_83 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c83
*+ bl_0_83 br_0_83 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c83
*+ bl_0_83 br_0_83 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c83
*+ bl_0_83 br_0_83 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c83
*+ bl_0_83 br_0_83 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c83
*+ bl_0_83 br_0_83 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c83
*+ bl_0_83 br_0_83 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c83
*+ bl_0_83 br_0_83 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c83
*+ bl_0_83 br_0_83 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c83
*+ bl_0_83 br_0_83 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c83
*+ bl_0_83 br_0_83 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c83
*+ bl_0_83 br_0_83 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c83
+ bl_0_83 br_0_83 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c84
+ bl_0_84 br_0_84 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c84
*+ bl_0_84 br_0_84 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c84
*+ bl_0_84 br_0_84 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c84
*+ bl_0_84 br_0_84 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c84
*+ bl_0_84 br_0_84 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c84
*+ bl_0_84 br_0_84 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c84
*+ bl_0_84 br_0_84 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c84
*+ bl_0_84 br_0_84 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c84
*+ bl_0_84 br_0_84 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c84
*+ bl_0_84 br_0_84 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c84
*+ bl_0_84 br_0_84 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c84
*+ bl_0_84 br_0_84 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c84
*+ bl_0_84 br_0_84 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c84
*+ bl_0_84 br_0_84 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c84
*+ bl_0_84 br_0_84 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c84
*+ bl_0_84 br_0_84 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c84
*+ bl_0_84 br_0_84 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c84
*+ bl_0_84 br_0_84 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c84
*+ bl_0_84 br_0_84 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c84
*+ bl_0_84 br_0_84 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c84
*+ bl_0_84 br_0_84 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c84
*+ bl_0_84 br_0_84 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c84
*+ bl_0_84 br_0_84 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c84
*+ bl_0_84 br_0_84 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c84
*+ bl_0_84 br_0_84 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c84
*+ bl_0_84 br_0_84 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c84
*+ bl_0_84 br_0_84 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c84
*+ bl_0_84 br_0_84 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c84
*+ bl_0_84 br_0_84 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c84
*+ bl_0_84 br_0_84 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c84
*+ bl_0_84 br_0_84 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c84
*+ bl_0_84 br_0_84 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c84
*+ bl_0_84 br_0_84 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c84
*+ bl_0_84 br_0_84 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c84
*+ bl_0_84 br_0_84 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c84
*+ bl_0_84 br_0_84 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c84
*+ bl_0_84 br_0_84 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c84
*+ bl_0_84 br_0_84 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c84
*+ bl_0_84 br_0_84 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c84
*+ bl_0_84 br_0_84 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c84
*+ bl_0_84 br_0_84 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c84
*+ bl_0_84 br_0_84 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c84
*+ bl_0_84 br_0_84 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c84
*+ bl_0_84 br_0_84 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c84
*+ bl_0_84 br_0_84 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c84
*+ bl_0_84 br_0_84 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c84
*+ bl_0_84 br_0_84 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c84
*+ bl_0_84 br_0_84 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c84
*+ bl_0_84 br_0_84 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c84
*+ bl_0_84 br_0_84 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c84
*+ bl_0_84 br_0_84 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c84
*+ bl_0_84 br_0_84 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c84
*+ bl_0_84 br_0_84 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c84
*+ bl_0_84 br_0_84 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c84
*+ bl_0_84 br_0_84 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c84
*+ bl_0_84 br_0_84 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c84
*+ bl_0_84 br_0_84 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c84
*+ bl_0_84 br_0_84 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c84
*+ bl_0_84 br_0_84 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c84
*+ bl_0_84 br_0_84 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c84
*+ bl_0_84 br_0_84 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c84
*+ bl_0_84 br_0_84 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c84
*+ bl_0_84 br_0_84 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c84
*+ bl_0_84 br_0_84 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c84
*+ bl_0_84 br_0_84 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c84
*+ bl_0_84 br_0_84 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c84
*+ bl_0_84 br_0_84 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c84
*+ bl_0_84 br_0_84 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c84
*+ bl_0_84 br_0_84 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c84
*+ bl_0_84 br_0_84 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c84
*+ bl_0_84 br_0_84 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c84
*+ bl_0_84 br_0_84 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c84
*+ bl_0_84 br_0_84 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c84
*+ bl_0_84 br_0_84 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c84
*+ bl_0_84 br_0_84 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c84
*+ bl_0_84 br_0_84 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c84
*+ bl_0_84 br_0_84 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c84
*+ bl_0_84 br_0_84 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c84
*+ bl_0_84 br_0_84 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c84
*+ bl_0_84 br_0_84 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c84
*+ bl_0_84 br_0_84 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c84
*+ bl_0_84 br_0_84 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c84
*+ bl_0_84 br_0_84 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c84
*+ bl_0_84 br_0_84 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c84
*+ bl_0_84 br_0_84 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c84
*+ bl_0_84 br_0_84 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c84
*+ bl_0_84 br_0_84 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c84
*+ bl_0_84 br_0_84 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c84
*+ bl_0_84 br_0_84 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c84
*+ bl_0_84 br_0_84 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c84
*+ bl_0_84 br_0_84 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c84
*+ bl_0_84 br_0_84 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c84
*+ bl_0_84 br_0_84 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c84
*+ bl_0_84 br_0_84 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c84
*+ bl_0_84 br_0_84 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c84
*+ bl_0_84 br_0_84 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c84
*+ bl_0_84 br_0_84 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c84
*+ bl_0_84 br_0_84 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c84
*+ bl_0_84 br_0_84 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c84
*+ bl_0_84 br_0_84 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c84
*+ bl_0_84 br_0_84 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c84
*+ bl_0_84 br_0_84 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c84
*+ bl_0_84 br_0_84 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c84
*+ bl_0_84 br_0_84 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c84
*+ bl_0_84 br_0_84 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c84
*+ bl_0_84 br_0_84 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c84
*+ bl_0_84 br_0_84 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c84
*+ bl_0_84 br_0_84 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c84
*+ bl_0_84 br_0_84 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c84
*+ bl_0_84 br_0_84 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c84
*+ bl_0_84 br_0_84 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c84
*+ bl_0_84 br_0_84 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c84
*+ bl_0_84 br_0_84 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c84
*+ bl_0_84 br_0_84 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c84
*+ bl_0_84 br_0_84 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c84
*+ bl_0_84 br_0_84 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c84
*+ bl_0_84 br_0_84 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c84
*+ bl_0_84 br_0_84 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c84
*+ bl_0_84 br_0_84 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c84
*+ bl_0_84 br_0_84 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c84
*+ bl_0_84 br_0_84 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c84
*+ bl_0_84 br_0_84 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c84
*+ bl_0_84 br_0_84 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c84
*+ bl_0_84 br_0_84 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c84
*+ bl_0_84 br_0_84 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c84
*+ bl_0_84 br_0_84 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c84
*+ bl_0_84 br_0_84 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c84
+ bl_0_84 br_0_84 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c85
+ bl_0_85 br_0_85 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c85
*+ bl_0_85 br_0_85 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c85
*+ bl_0_85 br_0_85 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c85
*+ bl_0_85 br_0_85 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c85
*+ bl_0_85 br_0_85 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c85
*+ bl_0_85 br_0_85 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c85
*+ bl_0_85 br_0_85 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c85
*+ bl_0_85 br_0_85 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c85
*+ bl_0_85 br_0_85 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c85
*+ bl_0_85 br_0_85 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c85
*+ bl_0_85 br_0_85 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c85
*+ bl_0_85 br_0_85 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c85
*+ bl_0_85 br_0_85 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c85
*+ bl_0_85 br_0_85 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c85
*+ bl_0_85 br_0_85 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c85
*+ bl_0_85 br_0_85 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c85
*+ bl_0_85 br_0_85 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c85
*+ bl_0_85 br_0_85 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c85
*+ bl_0_85 br_0_85 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c85
*+ bl_0_85 br_0_85 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c85
*+ bl_0_85 br_0_85 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c85
*+ bl_0_85 br_0_85 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c85
*+ bl_0_85 br_0_85 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c85
*+ bl_0_85 br_0_85 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c85
*+ bl_0_85 br_0_85 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c85
*+ bl_0_85 br_0_85 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c85
*+ bl_0_85 br_0_85 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c85
*+ bl_0_85 br_0_85 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c85
*+ bl_0_85 br_0_85 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c85
*+ bl_0_85 br_0_85 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c85
*+ bl_0_85 br_0_85 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c85
*+ bl_0_85 br_0_85 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c85
*+ bl_0_85 br_0_85 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c85
*+ bl_0_85 br_0_85 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c85
*+ bl_0_85 br_0_85 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c85
*+ bl_0_85 br_0_85 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c85
*+ bl_0_85 br_0_85 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c85
*+ bl_0_85 br_0_85 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c85
*+ bl_0_85 br_0_85 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c85
*+ bl_0_85 br_0_85 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c85
*+ bl_0_85 br_0_85 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c85
*+ bl_0_85 br_0_85 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c85
*+ bl_0_85 br_0_85 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c85
*+ bl_0_85 br_0_85 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c85
*+ bl_0_85 br_0_85 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c85
*+ bl_0_85 br_0_85 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c85
*+ bl_0_85 br_0_85 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c85
*+ bl_0_85 br_0_85 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c85
*+ bl_0_85 br_0_85 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c85
*+ bl_0_85 br_0_85 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c85
*+ bl_0_85 br_0_85 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c85
*+ bl_0_85 br_0_85 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c85
*+ bl_0_85 br_0_85 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c85
*+ bl_0_85 br_0_85 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c85
*+ bl_0_85 br_0_85 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c85
*+ bl_0_85 br_0_85 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c85
*+ bl_0_85 br_0_85 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c85
*+ bl_0_85 br_0_85 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c85
*+ bl_0_85 br_0_85 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c85
*+ bl_0_85 br_0_85 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c85
*+ bl_0_85 br_0_85 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c85
*+ bl_0_85 br_0_85 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c85
*+ bl_0_85 br_0_85 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c85
*+ bl_0_85 br_0_85 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c85
*+ bl_0_85 br_0_85 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c85
*+ bl_0_85 br_0_85 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c85
*+ bl_0_85 br_0_85 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c85
*+ bl_0_85 br_0_85 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c85
*+ bl_0_85 br_0_85 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c85
*+ bl_0_85 br_0_85 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c85
*+ bl_0_85 br_0_85 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c85
*+ bl_0_85 br_0_85 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c85
*+ bl_0_85 br_0_85 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c85
*+ bl_0_85 br_0_85 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c85
*+ bl_0_85 br_0_85 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c85
*+ bl_0_85 br_0_85 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c85
*+ bl_0_85 br_0_85 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c85
*+ bl_0_85 br_0_85 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c85
*+ bl_0_85 br_0_85 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c85
*+ bl_0_85 br_0_85 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c85
*+ bl_0_85 br_0_85 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c85
*+ bl_0_85 br_0_85 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c85
*+ bl_0_85 br_0_85 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c85
*+ bl_0_85 br_0_85 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c85
*+ bl_0_85 br_0_85 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c85
*+ bl_0_85 br_0_85 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c85
*+ bl_0_85 br_0_85 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c85
*+ bl_0_85 br_0_85 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c85
*+ bl_0_85 br_0_85 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c85
*+ bl_0_85 br_0_85 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c85
*+ bl_0_85 br_0_85 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c85
*+ bl_0_85 br_0_85 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c85
*+ bl_0_85 br_0_85 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c85
*+ bl_0_85 br_0_85 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c85
*+ bl_0_85 br_0_85 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c85
*+ bl_0_85 br_0_85 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c85
*+ bl_0_85 br_0_85 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c85
*+ bl_0_85 br_0_85 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c85
*+ bl_0_85 br_0_85 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c85
*+ bl_0_85 br_0_85 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c85
*+ bl_0_85 br_0_85 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c85
*+ bl_0_85 br_0_85 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c85
*+ bl_0_85 br_0_85 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c85
*+ bl_0_85 br_0_85 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c85
*+ bl_0_85 br_0_85 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c85
*+ bl_0_85 br_0_85 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c85
*+ bl_0_85 br_0_85 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c85
*+ bl_0_85 br_0_85 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c85
*+ bl_0_85 br_0_85 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c85
*+ bl_0_85 br_0_85 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c85
*+ bl_0_85 br_0_85 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c85
*+ bl_0_85 br_0_85 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c85
*+ bl_0_85 br_0_85 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c85
*+ bl_0_85 br_0_85 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c85
*+ bl_0_85 br_0_85 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c85
*+ bl_0_85 br_0_85 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c85
*+ bl_0_85 br_0_85 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c85
*+ bl_0_85 br_0_85 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c85
*+ bl_0_85 br_0_85 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c85
*+ bl_0_85 br_0_85 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c85
*+ bl_0_85 br_0_85 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c85
*+ bl_0_85 br_0_85 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c85
*+ bl_0_85 br_0_85 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c85
*+ bl_0_85 br_0_85 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c85
*+ bl_0_85 br_0_85 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c85
*+ bl_0_85 br_0_85 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c85
*+ bl_0_85 br_0_85 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c85
+ bl_0_85 br_0_85 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c86
+ bl_0_86 br_0_86 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c86
*+ bl_0_86 br_0_86 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c86
*+ bl_0_86 br_0_86 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c86
*+ bl_0_86 br_0_86 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c86
*+ bl_0_86 br_0_86 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c86
*+ bl_0_86 br_0_86 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c86
*+ bl_0_86 br_0_86 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c86
*+ bl_0_86 br_0_86 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c86
*+ bl_0_86 br_0_86 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c86
*+ bl_0_86 br_0_86 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c86
*+ bl_0_86 br_0_86 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c86
*+ bl_0_86 br_0_86 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c86
*+ bl_0_86 br_0_86 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c86
*+ bl_0_86 br_0_86 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c86
*+ bl_0_86 br_0_86 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c86
*+ bl_0_86 br_0_86 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c86
*+ bl_0_86 br_0_86 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c86
*+ bl_0_86 br_0_86 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c86
*+ bl_0_86 br_0_86 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c86
*+ bl_0_86 br_0_86 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c86
*+ bl_0_86 br_0_86 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c86
*+ bl_0_86 br_0_86 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c86
*+ bl_0_86 br_0_86 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c86
*+ bl_0_86 br_0_86 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c86
*+ bl_0_86 br_0_86 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c86
*+ bl_0_86 br_0_86 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c86
*+ bl_0_86 br_0_86 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c86
*+ bl_0_86 br_0_86 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c86
*+ bl_0_86 br_0_86 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c86
*+ bl_0_86 br_0_86 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c86
*+ bl_0_86 br_0_86 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c86
*+ bl_0_86 br_0_86 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c86
*+ bl_0_86 br_0_86 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c86
*+ bl_0_86 br_0_86 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c86
*+ bl_0_86 br_0_86 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c86
*+ bl_0_86 br_0_86 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c86
*+ bl_0_86 br_0_86 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c86
*+ bl_0_86 br_0_86 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c86
*+ bl_0_86 br_0_86 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c86
*+ bl_0_86 br_0_86 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c86
*+ bl_0_86 br_0_86 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c86
*+ bl_0_86 br_0_86 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c86
*+ bl_0_86 br_0_86 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c86
*+ bl_0_86 br_0_86 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c86
*+ bl_0_86 br_0_86 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c86
*+ bl_0_86 br_0_86 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c86
*+ bl_0_86 br_0_86 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c86
*+ bl_0_86 br_0_86 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c86
*+ bl_0_86 br_0_86 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c86
*+ bl_0_86 br_0_86 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c86
*+ bl_0_86 br_0_86 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c86
*+ bl_0_86 br_0_86 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c86
*+ bl_0_86 br_0_86 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c86
*+ bl_0_86 br_0_86 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c86
*+ bl_0_86 br_0_86 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c86
*+ bl_0_86 br_0_86 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c86
*+ bl_0_86 br_0_86 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c86
*+ bl_0_86 br_0_86 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c86
*+ bl_0_86 br_0_86 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c86
*+ bl_0_86 br_0_86 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c86
*+ bl_0_86 br_0_86 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c86
*+ bl_0_86 br_0_86 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c86
*+ bl_0_86 br_0_86 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c86
*+ bl_0_86 br_0_86 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c86
*+ bl_0_86 br_0_86 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c86
*+ bl_0_86 br_0_86 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c86
*+ bl_0_86 br_0_86 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c86
*+ bl_0_86 br_0_86 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c86
*+ bl_0_86 br_0_86 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c86
*+ bl_0_86 br_0_86 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c86
*+ bl_0_86 br_0_86 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c86
*+ bl_0_86 br_0_86 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c86
*+ bl_0_86 br_0_86 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c86
*+ bl_0_86 br_0_86 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c86
*+ bl_0_86 br_0_86 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c86
*+ bl_0_86 br_0_86 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c86
*+ bl_0_86 br_0_86 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c86
*+ bl_0_86 br_0_86 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c86
*+ bl_0_86 br_0_86 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c86
*+ bl_0_86 br_0_86 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c86
*+ bl_0_86 br_0_86 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c86
*+ bl_0_86 br_0_86 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c86
*+ bl_0_86 br_0_86 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c86
*+ bl_0_86 br_0_86 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c86
*+ bl_0_86 br_0_86 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c86
*+ bl_0_86 br_0_86 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c86
*+ bl_0_86 br_0_86 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c86
*+ bl_0_86 br_0_86 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c86
*+ bl_0_86 br_0_86 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c86
*+ bl_0_86 br_0_86 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c86
*+ bl_0_86 br_0_86 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c86
*+ bl_0_86 br_0_86 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c86
*+ bl_0_86 br_0_86 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c86
*+ bl_0_86 br_0_86 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c86
*+ bl_0_86 br_0_86 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c86
*+ bl_0_86 br_0_86 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c86
*+ bl_0_86 br_0_86 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c86
*+ bl_0_86 br_0_86 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c86
*+ bl_0_86 br_0_86 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c86
*+ bl_0_86 br_0_86 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c86
*+ bl_0_86 br_0_86 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c86
*+ bl_0_86 br_0_86 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c86
*+ bl_0_86 br_0_86 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c86
*+ bl_0_86 br_0_86 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c86
*+ bl_0_86 br_0_86 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c86
*+ bl_0_86 br_0_86 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c86
*+ bl_0_86 br_0_86 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c86
*+ bl_0_86 br_0_86 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c86
*+ bl_0_86 br_0_86 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c86
*+ bl_0_86 br_0_86 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c86
*+ bl_0_86 br_0_86 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c86
*+ bl_0_86 br_0_86 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c86
*+ bl_0_86 br_0_86 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c86
*+ bl_0_86 br_0_86 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c86
*+ bl_0_86 br_0_86 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c86
*+ bl_0_86 br_0_86 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c86
*+ bl_0_86 br_0_86 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c86
*+ bl_0_86 br_0_86 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c86
*+ bl_0_86 br_0_86 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c86
*+ bl_0_86 br_0_86 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c86
*+ bl_0_86 br_0_86 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c86
*+ bl_0_86 br_0_86 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c86
*+ bl_0_86 br_0_86 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c86
*+ bl_0_86 br_0_86 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c86
*+ bl_0_86 br_0_86 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c86
*+ bl_0_86 br_0_86 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c86
*+ bl_0_86 br_0_86 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c86
+ bl_0_86 br_0_86 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c87
+ bl_0_87 br_0_87 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c87
*+ bl_0_87 br_0_87 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c87
*+ bl_0_87 br_0_87 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c87
*+ bl_0_87 br_0_87 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c87
*+ bl_0_87 br_0_87 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c87
*+ bl_0_87 br_0_87 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c87
*+ bl_0_87 br_0_87 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c87
*+ bl_0_87 br_0_87 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c87
*+ bl_0_87 br_0_87 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c87
*+ bl_0_87 br_0_87 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c87
*+ bl_0_87 br_0_87 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c87
*+ bl_0_87 br_0_87 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c87
*+ bl_0_87 br_0_87 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c87
*+ bl_0_87 br_0_87 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c87
*+ bl_0_87 br_0_87 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c87
*+ bl_0_87 br_0_87 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c87
*+ bl_0_87 br_0_87 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c87
*+ bl_0_87 br_0_87 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c87
*+ bl_0_87 br_0_87 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c87
*+ bl_0_87 br_0_87 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c87
*+ bl_0_87 br_0_87 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c87
*+ bl_0_87 br_0_87 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c87
*+ bl_0_87 br_0_87 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c87
*+ bl_0_87 br_0_87 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c87
*+ bl_0_87 br_0_87 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c87
*+ bl_0_87 br_0_87 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c87
*+ bl_0_87 br_0_87 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c87
*+ bl_0_87 br_0_87 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c87
*+ bl_0_87 br_0_87 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c87
*+ bl_0_87 br_0_87 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c87
*+ bl_0_87 br_0_87 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c87
*+ bl_0_87 br_0_87 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c87
*+ bl_0_87 br_0_87 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c87
*+ bl_0_87 br_0_87 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c87
*+ bl_0_87 br_0_87 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c87
*+ bl_0_87 br_0_87 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c87
*+ bl_0_87 br_0_87 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c87
*+ bl_0_87 br_0_87 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c87
*+ bl_0_87 br_0_87 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c87
*+ bl_0_87 br_0_87 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c87
*+ bl_0_87 br_0_87 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c87
*+ bl_0_87 br_0_87 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c87
*+ bl_0_87 br_0_87 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c87
*+ bl_0_87 br_0_87 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c87
*+ bl_0_87 br_0_87 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c87
*+ bl_0_87 br_0_87 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c87
*+ bl_0_87 br_0_87 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c87
*+ bl_0_87 br_0_87 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c87
*+ bl_0_87 br_0_87 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c87
*+ bl_0_87 br_0_87 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c87
*+ bl_0_87 br_0_87 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c87
*+ bl_0_87 br_0_87 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c87
*+ bl_0_87 br_0_87 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c87
*+ bl_0_87 br_0_87 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c87
*+ bl_0_87 br_0_87 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c87
*+ bl_0_87 br_0_87 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c87
*+ bl_0_87 br_0_87 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c87
*+ bl_0_87 br_0_87 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c87
*+ bl_0_87 br_0_87 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c87
*+ bl_0_87 br_0_87 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c87
*+ bl_0_87 br_0_87 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c87
*+ bl_0_87 br_0_87 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c87
*+ bl_0_87 br_0_87 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c87
*+ bl_0_87 br_0_87 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c87
*+ bl_0_87 br_0_87 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c87
*+ bl_0_87 br_0_87 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c87
*+ bl_0_87 br_0_87 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c87
*+ bl_0_87 br_0_87 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c87
*+ bl_0_87 br_0_87 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c87
*+ bl_0_87 br_0_87 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c87
*+ bl_0_87 br_0_87 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c87
*+ bl_0_87 br_0_87 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c87
*+ bl_0_87 br_0_87 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c87
*+ bl_0_87 br_0_87 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c87
*+ bl_0_87 br_0_87 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c87
*+ bl_0_87 br_0_87 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c87
*+ bl_0_87 br_0_87 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c87
*+ bl_0_87 br_0_87 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c87
*+ bl_0_87 br_0_87 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c87
*+ bl_0_87 br_0_87 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c87
*+ bl_0_87 br_0_87 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c87
*+ bl_0_87 br_0_87 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c87
*+ bl_0_87 br_0_87 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c87
*+ bl_0_87 br_0_87 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c87
*+ bl_0_87 br_0_87 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c87
*+ bl_0_87 br_0_87 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c87
*+ bl_0_87 br_0_87 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c87
*+ bl_0_87 br_0_87 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c87
*+ bl_0_87 br_0_87 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c87
*+ bl_0_87 br_0_87 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c87
*+ bl_0_87 br_0_87 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c87
*+ bl_0_87 br_0_87 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c87
*+ bl_0_87 br_0_87 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c87
*+ bl_0_87 br_0_87 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c87
*+ bl_0_87 br_0_87 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c87
*+ bl_0_87 br_0_87 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c87
*+ bl_0_87 br_0_87 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c87
*+ bl_0_87 br_0_87 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c87
*+ bl_0_87 br_0_87 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c87
*+ bl_0_87 br_0_87 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c87
*+ bl_0_87 br_0_87 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c87
*+ bl_0_87 br_0_87 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c87
*+ bl_0_87 br_0_87 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c87
*+ bl_0_87 br_0_87 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c87
*+ bl_0_87 br_0_87 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c87
*+ bl_0_87 br_0_87 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c87
*+ bl_0_87 br_0_87 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c87
*+ bl_0_87 br_0_87 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c87
*+ bl_0_87 br_0_87 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c87
*+ bl_0_87 br_0_87 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c87
*+ bl_0_87 br_0_87 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c87
*+ bl_0_87 br_0_87 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c87
*+ bl_0_87 br_0_87 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c87
*+ bl_0_87 br_0_87 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c87
*+ bl_0_87 br_0_87 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c87
*+ bl_0_87 br_0_87 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c87
*+ bl_0_87 br_0_87 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c87
*+ bl_0_87 br_0_87 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c87
*+ bl_0_87 br_0_87 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c87
*+ bl_0_87 br_0_87 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c87
*+ bl_0_87 br_0_87 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c87
*+ bl_0_87 br_0_87 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c87
*+ bl_0_87 br_0_87 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c87
*+ bl_0_87 br_0_87 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c87
*+ bl_0_87 br_0_87 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c87
*+ bl_0_87 br_0_87 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c87
*+ bl_0_87 br_0_87 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c87
+ bl_0_87 br_0_87 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c88
+ bl_0_88 br_0_88 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c88
*+ bl_0_88 br_0_88 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c88
*+ bl_0_88 br_0_88 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c88
*+ bl_0_88 br_0_88 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c88
*+ bl_0_88 br_0_88 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c88
*+ bl_0_88 br_0_88 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c88
*+ bl_0_88 br_0_88 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c88
*+ bl_0_88 br_0_88 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c88
*+ bl_0_88 br_0_88 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c88
*+ bl_0_88 br_0_88 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c88
*+ bl_0_88 br_0_88 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c88
*+ bl_0_88 br_0_88 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c88
*+ bl_0_88 br_0_88 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c88
*+ bl_0_88 br_0_88 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c88
*+ bl_0_88 br_0_88 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c88
*+ bl_0_88 br_0_88 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c88
*+ bl_0_88 br_0_88 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c88
*+ bl_0_88 br_0_88 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c88
*+ bl_0_88 br_0_88 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c88
*+ bl_0_88 br_0_88 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c88
*+ bl_0_88 br_0_88 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c88
*+ bl_0_88 br_0_88 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c88
*+ bl_0_88 br_0_88 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c88
*+ bl_0_88 br_0_88 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c88
*+ bl_0_88 br_0_88 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c88
*+ bl_0_88 br_0_88 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c88
*+ bl_0_88 br_0_88 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c88
*+ bl_0_88 br_0_88 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c88
*+ bl_0_88 br_0_88 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c88
*+ bl_0_88 br_0_88 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c88
*+ bl_0_88 br_0_88 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c88
*+ bl_0_88 br_0_88 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c88
*+ bl_0_88 br_0_88 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c88
*+ bl_0_88 br_0_88 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c88
*+ bl_0_88 br_0_88 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c88
*+ bl_0_88 br_0_88 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c88
*+ bl_0_88 br_0_88 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c88
*+ bl_0_88 br_0_88 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c88
*+ bl_0_88 br_0_88 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c88
*+ bl_0_88 br_0_88 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c88
*+ bl_0_88 br_0_88 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c88
*+ bl_0_88 br_0_88 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c88
*+ bl_0_88 br_0_88 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c88
*+ bl_0_88 br_0_88 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c88
*+ bl_0_88 br_0_88 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c88
*+ bl_0_88 br_0_88 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c88
*+ bl_0_88 br_0_88 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c88
*+ bl_0_88 br_0_88 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c88
*+ bl_0_88 br_0_88 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c88
*+ bl_0_88 br_0_88 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c88
*+ bl_0_88 br_0_88 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c88
*+ bl_0_88 br_0_88 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c88
*+ bl_0_88 br_0_88 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c88
*+ bl_0_88 br_0_88 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c88
*+ bl_0_88 br_0_88 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c88
*+ bl_0_88 br_0_88 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c88
*+ bl_0_88 br_0_88 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c88
*+ bl_0_88 br_0_88 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c88
*+ bl_0_88 br_0_88 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c88
*+ bl_0_88 br_0_88 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c88
*+ bl_0_88 br_0_88 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c88
*+ bl_0_88 br_0_88 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c88
*+ bl_0_88 br_0_88 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c88
*+ bl_0_88 br_0_88 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c88
*+ bl_0_88 br_0_88 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c88
*+ bl_0_88 br_0_88 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c88
*+ bl_0_88 br_0_88 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c88
*+ bl_0_88 br_0_88 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c88
*+ bl_0_88 br_0_88 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c88
*+ bl_0_88 br_0_88 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c88
*+ bl_0_88 br_0_88 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c88
*+ bl_0_88 br_0_88 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c88
*+ bl_0_88 br_0_88 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c88
*+ bl_0_88 br_0_88 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c88
*+ bl_0_88 br_0_88 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c88
*+ bl_0_88 br_0_88 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c88
*+ bl_0_88 br_0_88 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c88
*+ bl_0_88 br_0_88 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c88
*+ bl_0_88 br_0_88 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c88
*+ bl_0_88 br_0_88 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c88
*+ bl_0_88 br_0_88 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c88
*+ bl_0_88 br_0_88 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c88
*+ bl_0_88 br_0_88 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c88
*+ bl_0_88 br_0_88 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c88
*+ bl_0_88 br_0_88 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c88
*+ bl_0_88 br_0_88 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c88
*+ bl_0_88 br_0_88 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c88
*+ bl_0_88 br_0_88 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c88
*+ bl_0_88 br_0_88 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c88
*+ bl_0_88 br_0_88 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c88
*+ bl_0_88 br_0_88 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c88
*+ bl_0_88 br_0_88 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c88
*+ bl_0_88 br_0_88 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c88
*+ bl_0_88 br_0_88 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c88
*+ bl_0_88 br_0_88 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c88
*+ bl_0_88 br_0_88 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c88
*+ bl_0_88 br_0_88 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c88
*+ bl_0_88 br_0_88 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c88
*+ bl_0_88 br_0_88 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c88
*+ bl_0_88 br_0_88 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c88
*+ bl_0_88 br_0_88 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c88
*+ bl_0_88 br_0_88 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c88
*+ bl_0_88 br_0_88 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c88
*+ bl_0_88 br_0_88 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c88
*+ bl_0_88 br_0_88 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c88
*+ bl_0_88 br_0_88 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c88
*+ bl_0_88 br_0_88 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c88
*+ bl_0_88 br_0_88 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c88
*+ bl_0_88 br_0_88 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c88
*+ bl_0_88 br_0_88 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c88
*+ bl_0_88 br_0_88 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c88
*+ bl_0_88 br_0_88 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c88
*+ bl_0_88 br_0_88 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c88
*+ bl_0_88 br_0_88 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c88
*+ bl_0_88 br_0_88 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c88
*+ bl_0_88 br_0_88 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c88
*+ bl_0_88 br_0_88 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c88
*+ bl_0_88 br_0_88 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c88
*+ bl_0_88 br_0_88 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c88
*+ bl_0_88 br_0_88 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c88
*+ bl_0_88 br_0_88 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c88
*+ bl_0_88 br_0_88 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c88
*+ bl_0_88 br_0_88 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c88
*+ bl_0_88 br_0_88 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c88
*+ bl_0_88 br_0_88 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c88
*+ bl_0_88 br_0_88 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c88
*+ bl_0_88 br_0_88 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c88
+ bl_0_88 br_0_88 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c89
+ bl_0_89 br_0_89 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c89
*+ bl_0_89 br_0_89 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c89
*+ bl_0_89 br_0_89 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c89
*+ bl_0_89 br_0_89 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c89
*+ bl_0_89 br_0_89 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c89
*+ bl_0_89 br_0_89 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c89
*+ bl_0_89 br_0_89 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c89
*+ bl_0_89 br_0_89 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c89
*+ bl_0_89 br_0_89 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c89
*+ bl_0_89 br_0_89 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c89
*+ bl_0_89 br_0_89 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c89
*+ bl_0_89 br_0_89 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c89
*+ bl_0_89 br_0_89 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c89
*+ bl_0_89 br_0_89 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c89
*+ bl_0_89 br_0_89 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c89
*+ bl_0_89 br_0_89 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c89
*+ bl_0_89 br_0_89 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c89
*+ bl_0_89 br_0_89 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c89
*+ bl_0_89 br_0_89 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c89
*+ bl_0_89 br_0_89 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c89
*+ bl_0_89 br_0_89 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c89
*+ bl_0_89 br_0_89 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c89
*+ bl_0_89 br_0_89 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c89
*+ bl_0_89 br_0_89 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c89
*+ bl_0_89 br_0_89 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c89
*+ bl_0_89 br_0_89 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c89
*+ bl_0_89 br_0_89 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c89
*+ bl_0_89 br_0_89 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c89
*+ bl_0_89 br_0_89 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c89
*+ bl_0_89 br_0_89 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c89
*+ bl_0_89 br_0_89 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c89
*+ bl_0_89 br_0_89 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c89
*+ bl_0_89 br_0_89 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c89
*+ bl_0_89 br_0_89 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c89
*+ bl_0_89 br_0_89 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c89
*+ bl_0_89 br_0_89 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c89
*+ bl_0_89 br_0_89 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c89
*+ bl_0_89 br_0_89 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c89
*+ bl_0_89 br_0_89 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c89
*+ bl_0_89 br_0_89 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c89
*+ bl_0_89 br_0_89 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c89
*+ bl_0_89 br_0_89 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c89
*+ bl_0_89 br_0_89 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c89
*+ bl_0_89 br_0_89 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c89
*+ bl_0_89 br_0_89 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c89
*+ bl_0_89 br_0_89 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c89
*+ bl_0_89 br_0_89 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c89
*+ bl_0_89 br_0_89 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c89
*+ bl_0_89 br_0_89 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c89
*+ bl_0_89 br_0_89 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c89
*+ bl_0_89 br_0_89 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c89
*+ bl_0_89 br_0_89 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c89
*+ bl_0_89 br_0_89 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c89
*+ bl_0_89 br_0_89 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c89
*+ bl_0_89 br_0_89 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c89
*+ bl_0_89 br_0_89 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c89
*+ bl_0_89 br_0_89 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c89
*+ bl_0_89 br_0_89 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c89
*+ bl_0_89 br_0_89 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c89
*+ bl_0_89 br_0_89 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c89
*+ bl_0_89 br_0_89 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c89
*+ bl_0_89 br_0_89 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c89
*+ bl_0_89 br_0_89 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c89
*+ bl_0_89 br_0_89 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c89
*+ bl_0_89 br_0_89 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c89
*+ bl_0_89 br_0_89 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c89
*+ bl_0_89 br_0_89 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c89
*+ bl_0_89 br_0_89 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c89
*+ bl_0_89 br_0_89 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c89
*+ bl_0_89 br_0_89 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c89
*+ bl_0_89 br_0_89 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c89
*+ bl_0_89 br_0_89 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c89
*+ bl_0_89 br_0_89 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c89
*+ bl_0_89 br_0_89 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c89
*+ bl_0_89 br_0_89 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c89
*+ bl_0_89 br_0_89 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c89
*+ bl_0_89 br_0_89 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c89
*+ bl_0_89 br_0_89 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c89
*+ bl_0_89 br_0_89 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c89
*+ bl_0_89 br_0_89 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c89
*+ bl_0_89 br_0_89 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c89
*+ bl_0_89 br_0_89 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c89
*+ bl_0_89 br_0_89 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c89
*+ bl_0_89 br_0_89 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c89
*+ bl_0_89 br_0_89 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c89
*+ bl_0_89 br_0_89 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c89
*+ bl_0_89 br_0_89 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c89
*+ bl_0_89 br_0_89 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c89
*+ bl_0_89 br_0_89 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c89
*+ bl_0_89 br_0_89 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c89
*+ bl_0_89 br_0_89 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c89
*+ bl_0_89 br_0_89 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c89
*+ bl_0_89 br_0_89 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c89
*+ bl_0_89 br_0_89 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c89
*+ bl_0_89 br_0_89 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c89
*+ bl_0_89 br_0_89 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c89
*+ bl_0_89 br_0_89 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c89
*+ bl_0_89 br_0_89 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c89
*+ bl_0_89 br_0_89 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c89
*+ bl_0_89 br_0_89 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c89
*+ bl_0_89 br_0_89 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c89
*+ bl_0_89 br_0_89 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c89
*+ bl_0_89 br_0_89 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c89
*+ bl_0_89 br_0_89 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c89
*+ bl_0_89 br_0_89 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c89
*+ bl_0_89 br_0_89 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c89
*+ bl_0_89 br_0_89 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c89
*+ bl_0_89 br_0_89 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c89
*+ bl_0_89 br_0_89 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c89
*+ bl_0_89 br_0_89 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c89
*+ bl_0_89 br_0_89 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c89
*+ bl_0_89 br_0_89 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c89
*+ bl_0_89 br_0_89 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c89
*+ bl_0_89 br_0_89 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c89
*+ bl_0_89 br_0_89 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c89
*+ bl_0_89 br_0_89 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c89
*+ bl_0_89 br_0_89 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c89
*+ bl_0_89 br_0_89 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c89
*+ bl_0_89 br_0_89 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c89
*+ bl_0_89 br_0_89 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c89
*+ bl_0_89 br_0_89 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c89
*+ bl_0_89 br_0_89 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c89
*+ bl_0_89 br_0_89 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c89
*+ bl_0_89 br_0_89 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c89
*+ bl_0_89 br_0_89 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c89
*+ bl_0_89 br_0_89 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c89
*+ bl_0_89 br_0_89 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c89
+ bl_0_89 br_0_89 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c90
+ bl_0_90 br_0_90 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c90
*+ bl_0_90 br_0_90 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c90
*+ bl_0_90 br_0_90 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c90
*+ bl_0_90 br_0_90 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c90
*+ bl_0_90 br_0_90 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c90
*+ bl_0_90 br_0_90 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c90
*+ bl_0_90 br_0_90 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c90
*+ bl_0_90 br_0_90 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c90
*+ bl_0_90 br_0_90 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c90
*+ bl_0_90 br_0_90 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c90
*+ bl_0_90 br_0_90 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c90
*+ bl_0_90 br_0_90 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c90
*+ bl_0_90 br_0_90 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c90
*+ bl_0_90 br_0_90 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c90
*+ bl_0_90 br_0_90 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c90
*+ bl_0_90 br_0_90 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c90
*+ bl_0_90 br_0_90 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c90
*+ bl_0_90 br_0_90 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c90
*+ bl_0_90 br_0_90 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c90
*+ bl_0_90 br_0_90 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c90
*+ bl_0_90 br_0_90 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c90
*+ bl_0_90 br_0_90 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c90
*+ bl_0_90 br_0_90 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c90
*+ bl_0_90 br_0_90 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c90
*+ bl_0_90 br_0_90 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c90
*+ bl_0_90 br_0_90 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c90
*+ bl_0_90 br_0_90 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c90
*+ bl_0_90 br_0_90 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c90
*+ bl_0_90 br_0_90 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c90
*+ bl_0_90 br_0_90 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c90
*+ bl_0_90 br_0_90 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c90
*+ bl_0_90 br_0_90 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c90
*+ bl_0_90 br_0_90 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c90
*+ bl_0_90 br_0_90 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c90
*+ bl_0_90 br_0_90 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c90
*+ bl_0_90 br_0_90 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c90
*+ bl_0_90 br_0_90 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c90
*+ bl_0_90 br_0_90 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c90
*+ bl_0_90 br_0_90 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c90
*+ bl_0_90 br_0_90 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c90
*+ bl_0_90 br_0_90 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c90
*+ bl_0_90 br_0_90 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c90
*+ bl_0_90 br_0_90 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c90
*+ bl_0_90 br_0_90 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c90
*+ bl_0_90 br_0_90 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c90
*+ bl_0_90 br_0_90 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c90
*+ bl_0_90 br_0_90 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c90
*+ bl_0_90 br_0_90 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c90
*+ bl_0_90 br_0_90 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c90
*+ bl_0_90 br_0_90 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c90
*+ bl_0_90 br_0_90 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c90
*+ bl_0_90 br_0_90 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c90
*+ bl_0_90 br_0_90 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c90
*+ bl_0_90 br_0_90 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c90
*+ bl_0_90 br_0_90 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c90
*+ bl_0_90 br_0_90 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c90
*+ bl_0_90 br_0_90 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c90
*+ bl_0_90 br_0_90 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c90
*+ bl_0_90 br_0_90 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c90
*+ bl_0_90 br_0_90 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c90
*+ bl_0_90 br_0_90 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c90
*+ bl_0_90 br_0_90 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c90
*+ bl_0_90 br_0_90 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c90
*+ bl_0_90 br_0_90 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c90
*+ bl_0_90 br_0_90 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c90
*+ bl_0_90 br_0_90 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c90
*+ bl_0_90 br_0_90 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c90
*+ bl_0_90 br_0_90 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c90
*+ bl_0_90 br_0_90 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c90
*+ bl_0_90 br_0_90 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c90
*+ bl_0_90 br_0_90 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c90
*+ bl_0_90 br_0_90 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c90
*+ bl_0_90 br_0_90 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c90
*+ bl_0_90 br_0_90 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c90
*+ bl_0_90 br_0_90 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c90
*+ bl_0_90 br_0_90 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c90
*+ bl_0_90 br_0_90 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c90
*+ bl_0_90 br_0_90 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c90
*+ bl_0_90 br_0_90 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c90
*+ bl_0_90 br_0_90 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c90
*+ bl_0_90 br_0_90 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c90
*+ bl_0_90 br_0_90 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c90
*+ bl_0_90 br_0_90 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c90
*+ bl_0_90 br_0_90 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c90
*+ bl_0_90 br_0_90 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c90
*+ bl_0_90 br_0_90 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c90
*+ bl_0_90 br_0_90 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c90
*+ bl_0_90 br_0_90 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c90
*+ bl_0_90 br_0_90 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c90
*+ bl_0_90 br_0_90 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c90
*+ bl_0_90 br_0_90 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c90
*+ bl_0_90 br_0_90 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c90
*+ bl_0_90 br_0_90 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c90
*+ bl_0_90 br_0_90 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c90
*+ bl_0_90 br_0_90 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c90
*+ bl_0_90 br_0_90 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c90
*+ bl_0_90 br_0_90 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c90
*+ bl_0_90 br_0_90 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c90
*+ bl_0_90 br_0_90 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c90
*+ bl_0_90 br_0_90 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c90
*+ bl_0_90 br_0_90 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c90
*+ bl_0_90 br_0_90 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c90
*+ bl_0_90 br_0_90 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c90
*+ bl_0_90 br_0_90 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c90
*+ bl_0_90 br_0_90 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c90
*+ bl_0_90 br_0_90 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c90
*+ bl_0_90 br_0_90 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c90
*+ bl_0_90 br_0_90 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c90
*+ bl_0_90 br_0_90 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c90
*+ bl_0_90 br_0_90 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c90
*+ bl_0_90 br_0_90 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c90
*+ bl_0_90 br_0_90 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c90
*+ bl_0_90 br_0_90 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c90
*+ bl_0_90 br_0_90 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c90
*+ bl_0_90 br_0_90 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c90
*+ bl_0_90 br_0_90 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c90
*+ bl_0_90 br_0_90 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c90
*+ bl_0_90 br_0_90 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c90
*+ bl_0_90 br_0_90 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c90
*+ bl_0_90 br_0_90 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c90
*+ bl_0_90 br_0_90 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c90
*+ bl_0_90 br_0_90 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c90
*+ bl_0_90 br_0_90 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c90
*+ bl_0_90 br_0_90 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c90
*+ bl_0_90 br_0_90 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c90
*+ bl_0_90 br_0_90 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c90
*+ bl_0_90 br_0_90 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c90
+ bl_0_90 br_0_90 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c91
+ bl_0_91 br_0_91 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c91
*+ bl_0_91 br_0_91 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c91
*+ bl_0_91 br_0_91 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c91
*+ bl_0_91 br_0_91 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c91
*+ bl_0_91 br_0_91 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c91
*+ bl_0_91 br_0_91 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c91
*+ bl_0_91 br_0_91 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c91
*+ bl_0_91 br_0_91 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c91
*+ bl_0_91 br_0_91 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c91
*+ bl_0_91 br_0_91 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c91
*+ bl_0_91 br_0_91 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c91
*+ bl_0_91 br_0_91 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c91
*+ bl_0_91 br_0_91 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c91
*+ bl_0_91 br_0_91 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c91
*+ bl_0_91 br_0_91 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c91
*+ bl_0_91 br_0_91 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c91
*+ bl_0_91 br_0_91 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c91
*+ bl_0_91 br_0_91 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c91
*+ bl_0_91 br_0_91 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c91
*+ bl_0_91 br_0_91 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c91
*+ bl_0_91 br_0_91 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c91
*+ bl_0_91 br_0_91 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c91
*+ bl_0_91 br_0_91 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c91
*+ bl_0_91 br_0_91 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c91
*+ bl_0_91 br_0_91 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c91
*+ bl_0_91 br_0_91 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c91
*+ bl_0_91 br_0_91 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c91
*+ bl_0_91 br_0_91 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c91
*+ bl_0_91 br_0_91 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c91
*+ bl_0_91 br_0_91 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c91
*+ bl_0_91 br_0_91 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c91
*+ bl_0_91 br_0_91 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c91
*+ bl_0_91 br_0_91 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c91
*+ bl_0_91 br_0_91 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c91
*+ bl_0_91 br_0_91 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c91
*+ bl_0_91 br_0_91 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c91
*+ bl_0_91 br_0_91 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c91
*+ bl_0_91 br_0_91 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c91
*+ bl_0_91 br_0_91 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c91
*+ bl_0_91 br_0_91 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c91
*+ bl_0_91 br_0_91 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c91
*+ bl_0_91 br_0_91 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c91
*+ bl_0_91 br_0_91 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c91
*+ bl_0_91 br_0_91 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c91
*+ bl_0_91 br_0_91 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c91
*+ bl_0_91 br_0_91 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c91
*+ bl_0_91 br_0_91 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c91
*+ bl_0_91 br_0_91 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c91
*+ bl_0_91 br_0_91 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c91
*+ bl_0_91 br_0_91 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c91
*+ bl_0_91 br_0_91 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c91
*+ bl_0_91 br_0_91 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c91
*+ bl_0_91 br_0_91 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c91
*+ bl_0_91 br_0_91 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c91
*+ bl_0_91 br_0_91 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c91
*+ bl_0_91 br_0_91 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c91
*+ bl_0_91 br_0_91 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c91
*+ bl_0_91 br_0_91 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c91
*+ bl_0_91 br_0_91 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c91
*+ bl_0_91 br_0_91 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c91
*+ bl_0_91 br_0_91 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c91
*+ bl_0_91 br_0_91 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c91
*+ bl_0_91 br_0_91 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c91
*+ bl_0_91 br_0_91 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c91
*+ bl_0_91 br_0_91 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c91
*+ bl_0_91 br_0_91 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c91
*+ bl_0_91 br_0_91 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c91
*+ bl_0_91 br_0_91 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c91
*+ bl_0_91 br_0_91 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c91
*+ bl_0_91 br_0_91 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c91
*+ bl_0_91 br_0_91 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c91
*+ bl_0_91 br_0_91 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c91
*+ bl_0_91 br_0_91 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c91
*+ bl_0_91 br_0_91 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c91
*+ bl_0_91 br_0_91 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c91
*+ bl_0_91 br_0_91 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c91
*+ bl_0_91 br_0_91 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c91
*+ bl_0_91 br_0_91 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c91
*+ bl_0_91 br_0_91 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c91
*+ bl_0_91 br_0_91 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c91
*+ bl_0_91 br_0_91 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c91
*+ bl_0_91 br_0_91 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c91
*+ bl_0_91 br_0_91 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c91
*+ bl_0_91 br_0_91 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c91
*+ bl_0_91 br_0_91 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c91
*+ bl_0_91 br_0_91 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c91
*+ bl_0_91 br_0_91 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c91
*+ bl_0_91 br_0_91 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c91
*+ bl_0_91 br_0_91 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c91
*+ bl_0_91 br_0_91 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c91
*+ bl_0_91 br_0_91 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c91
*+ bl_0_91 br_0_91 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c91
*+ bl_0_91 br_0_91 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c91
*+ bl_0_91 br_0_91 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c91
*+ bl_0_91 br_0_91 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c91
*+ bl_0_91 br_0_91 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c91
*+ bl_0_91 br_0_91 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c91
*+ bl_0_91 br_0_91 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c91
*+ bl_0_91 br_0_91 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c91
*+ bl_0_91 br_0_91 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c91
*+ bl_0_91 br_0_91 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c91
*+ bl_0_91 br_0_91 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c91
*+ bl_0_91 br_0_91 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c91
*+ bl_0_91 br_0_91 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c91
*+ bl_0_91 br_0_91 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c91
*+ bl_0_91 br_0_91 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c91
*+ bl_0_91 br_0_91 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c91
*+ bl_0_91 br_0_91 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c91
*+ bl_0_91 br_0_91 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c91
*+ bl_0_91 br_0_91 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c91
*+ bl_0_91 br_0_91 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c91
*+ bl_0_91 br_0_91 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c91
*+ bl_0_91 br_0_91 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c91
*+ bl_0_91 br_0_91 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c91
*+ bl_0_91 br_0_91 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c91
*+ bl_0_91 br_0_91 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c91
*+ bl_0_91 br_0_91 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c91
*+ bl_0_91 br_0_91 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c91
*+ bl_0_91 br_0_91 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c91
*+ bl_0_91 br_0_91 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c91
*+ bl_0_91 br_0_91 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c91
*+ bl_0_91 br_0_91 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c91
*+ bl_0_91 br_0_91 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c91
*+ bl_0_91 br_0_91 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c91
*+ bl_0_91 br_0_91 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c91
*+ bl_0_91 br_0_91 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c91
*+ bl_0_91 br_0_91 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c91
+ bl_0_91 br_0_91 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c92
+ bl_0_92 br_0_92 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c92
*+ bl_0_92 br_0_92 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c92
*+ bl_0_92 br_0_92 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c92
*+ bl_0_92 br_0_92 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c92
*+ bl_0_92 br_0_92 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c92
*+ bl_0_92 br_0_92 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c92
*+ bl_0_92 br_0_92 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c92
*+ bl_0_92 br_0_92 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c92
*+ bl_0_92 br_0_92 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c92
*+ bl_0_92 br_0_92 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c92
*+ bl_0_92 br_0_92 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c92
*+ bl_0_92 br_0_92 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c92
*+ bl_0_92 br_0_92 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c92
*+ bl_0_92 br_0_92 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c92
*+ bl_0_92 br_0_92 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c92
*+ bl_0_92 br_0_92 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c92
*+ bl_0_92 br_0_92 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c92
*+ bl_0_92 br_0_92 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c92
*+ bl_0_92 br_0_92 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c92
*+ bl_0_92 br_0_92 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c92
*+ bl_0_92 br_0_92 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c92
*+ bl_0_92 br_0_92 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c92
*+ bl_0_92 br_0_92 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c92
*+ bl_0_92 br_0_92 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c92
*+ bl_0_92 br_0_92 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c92
*+ bl_0_92 br_0_92 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c92
*+ bl_0_92 br_0_92 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c92
*+ bl_0_92 br_0_92 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c92
*+ bl_0_92 br_0_92 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c92
*+ bl_0_92 br_0_92 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c92
*+ bl_0_92 br_0_92 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c92
*+ bl_0_92 br_0_92 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c92
*+ bl_0_92 br_0_92 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c92
*+ bl_0_92 br_0_92 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c92
*+ bl_0_92 br_0_92 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c92
*+ bl_0_92 br_0_92 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c92
*+ bl_0_92 br_0_92 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c92
*+ bl_0_92 br_0_92 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c92
*+ bl_0_92 br_0_92 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c92
*+ bl_0_92 br_0_92 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c92
*+ bl_0_92 br_0_92 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c92
*+ bl_0_92 br_0_92 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c92
*+ bl_0_92 br_0_92 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c92
*+ bl_0_92 br_0_92 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c92
*+ bl_0_92 br_0_92 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c92
*+ bl_0_92 br_0_92 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c92
*+ bl_0_92 br_0_92 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c92
*+ bl_0_92 br_0_92 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c92
*+ bl_0_92 br_0_92 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c92
*+ bl_0_92 br_0_92 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c92
*+ bl_0_92 br_0_92 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c92
*+ bl_0_92 br_0_92 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c92
*+ bl_0_92 br_0_92 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c92
*+ bl_0_92 br_0_92 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c92
*+ bl_0_92 br_0_92 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c92
*+ bl_0_92 br_0_92 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c92
*+ bl_0_92 br_0_92 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c92
*+ bl_0_92 br_0_92 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c92
*+ bl_0_92 br_0_92 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c92
*+ bl_0_92 br_0_92 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c92
*+ bl_0_92 br_0_92 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c92
*+ bl_0_92 br_0_92 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c92
*+ bl_0_92 br_0_92 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c92
*+ bl_0_92 br_0_92 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c92
*+ bl_0_92 br_0_92 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c92
*+ bl_0_92 br_0_92 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c92
*+ bl_0_92 br_0_92 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c92
*+ bl_0_92 br_0_92 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c92
*+ bl_0_92 br_0_92 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c92
*+ bl_0_92 br_0_92 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c92
*+ bl_0_92 br_0_92 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c92
*+ bl_0_92 br_0_92 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c92
*+ bl_0_92 br_0_92 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c92
*+ bl_0_92 br_0_92 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c92
*+ bl_0_92 br_0_92 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c92
*+ bl_0_92 br_0_92 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c92
*+ bl_0_92 br_0_92 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c92
*+ bl_0_92 br_0_92 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c92
*+ bl_0_92 br_0_92 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c92
*+ bl_0_92 br_0_92 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c92
*+ bl_0_92 br_0_92 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c92
*+ bl_0_92 br_0_92 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c92
*+ bl_0_92 br_0_92 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c92
*+ bl_0_92 br_0_92 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c92
*+ bl_0_92 br_0_92 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c92
*+ bl_0_92 br_0_92 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c92
*+ bl_0_92 br_0_92 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c92
*+ bl_0_92 br_0_92 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c92
*+ bl_0_92 br_0_92 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c92
*+ bl_0_92 br_0_92 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c92
*+ bl_0_92 br_0_92 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c92
*+ bl_0_92 br_0_92 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c92
*+ bl_0_92 br_0_92 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c92
*+ bl_0_92 br_0_92 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c92
*+ bl_0_92 br_0_92 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c92
*+ bl_0_92 br_0_92 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c92
*+ bl_0_92 br_0_92 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c92
*+ bl_0_92 br_0_92 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c92
*+ bl_0_92 br_0_92 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c92
*+ bl_0_92 br_0_92 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c92
*+ bl_0_92 br_0_92 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c92
*+ bl_0_92 br_0_92 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c92
*+ bl_0_92 br_0_92 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c92
*+ bl_0_92 br_0_92 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c92
*+ bl_0_92 br_0_92 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c92
*+ bl_0_92 br_0_92 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c92
*+ bl_0_92 br_0_92 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c92
*+ bl_0_92 br_0_92 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c92
*+ bl_0_92 br_0_92 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c92
*+ bl_0_92 br_0_92 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c92
*+ bl_0_92 br_0_92 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c92
*+ bl_0_92 br_0_92 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c92
*+ bl_0_92 br_0_92 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c92
*+ bl_0_92 br_0_92 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c92
*+ bl_0_92 br_0_92 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c92
*+ bl_0_92 br_0_92 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c92
*+ bl_0_92 br_0_92 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c92
*+ bl_0_92 br_0_92 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c92
*+ bl_0_92 br_0_92 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c92
*+ bl_0_92 br_0_92 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c92
*+ bl_0_92 br_0_92 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c92
*+ bl_0_92 br_0_92 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c92
*+ bl_0_92 br_0_92 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c92
*+ bl_0_92 br_0_92 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c92
*+ bl_0_92 br_0_92 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c92
*+ bl_0_92 br_0_92 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c92
*+ bl_0_92 br_0_92 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c92
+ bl_0_92 br_0_92 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c93
+ bl_0_93 br_0_93 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c93
*+ bl_0_93 br_0_93 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c93
*+ bl_0_93 br_0_93 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c93
*+ bl_0_93 br_0_93 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c93
*+ bl_0_93 br_0_93 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c93
*+ bl_0_93 br_0_93 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c93
*+ bl_0_93 br_0_93 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c93
*+ bl_0_93 br_0_93 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c93
*+ bl_0_93 br_0_93 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c93
*+ bl_0_93 br_0_93 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c93
*+ bl_0_93 br_0_93 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c93
*+ bl_0_93 br_0_93 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c93
*+ bl_0_93 br_0_93 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c93
*+ bl_0_93 br_0_93 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c93
*+ bl_0_93 br_0_93 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c93
*+ bl_0_93 br_0_93 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c93
*+ bl_0_93 br_0_93 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c93
*+ bl_0_93 br_0_93 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c93
*+ bl_0_93 br_0_93 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c93
*+ bl_0_93 br_0_93 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c93
*+ bl_0_93 br_0_93 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c93
*+ bl_0_93 br_0_93 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c93
*+ bl_0_93 br_0_93 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c93
*+ bl_0_93 br_0_93 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c93
*+ bl_0_93 br_0_93 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c93
*+ bl_0_93 br_0_93 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c93
*+ bl_0_93 br_0_93 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c93
*+ bl_0_93 br_0_93 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c93
*+ bl_0_93 br_0_93 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c93
*+ bl_0_93 br_0_93 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c93
*+ bl_0_93 br_0_93 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c93
*+ bl_0_93 br_0_93 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c93
*+ bl_0_93 br_0_93 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c93
*+ bl_0_93 br_0_93 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c93
*+ bl_0_93 br_0_93 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c93
*+ bl_0_93 br_0_93 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c93
*+ bl_0_93 br_0_93 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c93
*+ bl_0_93 br_0_93 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c93
*+ bl_0_93 br_0_93 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c93
*+ bl_0_93 br_0_93 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c93
*+ bl_0_93 br_0_93 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c93
*+ bl_0_93 br_0_93 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c93
*+ bl_0_93 br_0_93 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c93
*+ bl_0_93 br_0_93 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c93
*+ bl_0_93 br_0_93 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c93
*+ bl_0_93 br_0_93 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c93
*+ bl_0_93 br_0_93 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c93
*+ bl_0_93 br_0_93 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c93
*+ bl_0_93 br_0_93 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c93
*+ bl_0_93 br_0_93 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c93
*+ bl_0_93 br_0_93 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c93
*+ bl_0_93 br_0_93 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c93
*+ bl_0_93 br_0_93 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c93
*+ bl_0_93 br_0_93 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c93
*+ bl_0_93 br_0_93 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c93
*+ bl_0_93 br_0_93 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c93
*+ bl_0_93 br_0_93 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c93
*+ bl_0_93 br_0_93 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c93
*+ bl_0_93 br_0_93 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c93
*+ bl_0_93 br_0_93 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c93
*+ bl_0_93 br_0_93 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c93
*+ bl_0_93 br_0_93 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c93
*+ bl_0_93 br_0_93 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c93
*+ bl_0_93 br_0_93 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c93
*+ bl_0_93 br_0_93 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c93
*+ bl_0_93 br_0_93 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c93
*+ bl_0_93 br_0_93 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c93
*+ bl_0_93 br_0_93 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c93
*+ bl_0_93 br_0_93 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c93
*+ bl_0_93 br_0_93 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c93
*+ bl_0_93 br_0_93 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c93
*+ bl_0_93 br_0_93 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c93
*+ bl_0_93 br_0_93 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c93
*+ bl_0_93 br_0_93 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c93
*+ bl_0_93 br_0_93 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c93
*+ bl_0_93 br_0_93 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c93
*+ bl_0_93 br_0_93 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c93
*+ bl_0_93 br_0_93 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c93
*+ bl_0_93 br_0_93 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c93
*+ bl_0_93 br_0_93 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c93
*+ bl_0_93 br_0_93 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c93
*+ bl_0_93 br_0_93 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c93
*+ bl_0_93 br_0_93 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c93
*+ bl_0_93 br_0_93 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c93
*+ bl_0_93 br_0_93 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c93
*+ bl_0_93 br_0_93 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c93
*+ bl_0_93 br_0_93 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c93
*+ bl_0_93 br_0_93 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c93
*+ bl_0_93 br_0_93 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c93
*+ bl_0_93 br_0_93 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c93
*+ bl_0_93 br_0_93 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c93
*+ bl_0_93 br_0_93 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c93
*+ bl_0_93 br_0_93 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c93
*+ bl_0_93 br_0_93 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c93
*+ bl_0_93 br_0_93 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c93
*+ bl_0_93 br_0_93 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c93
*+ bl_0_93 br_0_93 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c93
*+ bl_0_93 br_0_93 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c93
*+ bl_0_93 br_0_93 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c93
*+ bl_0_93 br_0_93 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c93
*+ bl_0_93 br_0_93 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c93
*+ bl_0_93 br_0_93 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c93
*+ bl_0_93 br_0_93 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c93
*+ bl_0_93 br_0_93 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c93
*+ bl_0_93 br_0_93 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c93
*+ bl_0_93 br_0_93 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c93
*+ bl_0_93 br_0_93 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c93
*+ bl_0_93 br_0_93 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c93
*+ bl_0_93 br_0_93 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c93
*+ bl_0_93 br_0_93 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c93
*+ bl_0_93 br_0_93 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c93
*+ bl_0_93 br_0_93 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c93
*+ bl_0_93 br_0_93 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c93
*+ bl_0_93 br_0_93 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c93
*+ bl_0_93 br_0_93 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c93
*+ bl_0_93 br_0_93 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c93
*+ bl_0_93 br_0_93 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c93
*+ bl_0_93 br_0_93 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c93
*+ bl_0_93 br_0_93 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c93
*+ bl_0_93 br_0_93 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c93
*+ bl_0_93 br_0_93 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c93
*+ bl_0_93 br_0_93 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c93
*+ bl_0_93 br_0_93 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c93
*+ bl_0_93 br_0_93 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c93
*+ bl_0_93 br_0_93 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c93
*+ bl_0_93 br_0_93 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c93
*+ bl_0_93 br_0_93 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c93
+ bl_0_93 br_0_93 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c94
+ bl_0_94 br_0_94 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c94
*+ bl_0_94 br_0_94 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c94
*+ bl_0_94 br_0_94 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c94
*+ bl_0_94 br_0_94 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c94
*+ bl_0_94 br_0_94 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c94
*+ bl_0_94 br_0_94 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c94
*+ bl_0_94 br_0_94 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c94
*+ bl_0_94 br_0_94 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c94
*+ bl_0_94 br_0_94 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c94
*+ bl_0_94 br_0_94 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c94
*+ bl_0_94 br_0_94 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c94
*+ bl_0_94 br_0_94 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c94
*+ bl_0_94 br_0_94 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c94
*+ bl_0_94 br_0_94 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c94
*+ bl_0_94 br_0_94 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c94
*+ bl_0_94 br_0_94 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c94
*+ bl_0_94 br_0_94 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c94
*+ bl_0_94 br_0_94 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c94
*+ bl_0_94 br_0_94 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c94
*+ bl_0_94 br_0_94 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c94
*+ bl_0_94 br_0_94 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c94
*+ bl_0_94 br_0_94 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c94
*+ bl_0_94 br_0_94 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c94
*+ bl_0_94 br_0_94 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c94
*+ bl_0_94 br_0_94 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c94
*+ bl_0_94 br_0_94 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c94
*+ bl_0_94 br_0_94 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c94
*+ bl_0_94 br_0_94 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c94
*+ bl_0_94 br_0_94 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c94
*+ bl_0_94 br_0_94 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c94
*+ bl_0_94 br_0_94 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c94
*+ bl_0_94 br_0_94 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c94
*+ bl_0_94 br_0_94 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c94
*+ bl_0_94 br_0_94 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c94
*+ bl_0_94 br_0_94 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c94
*+ bl_0_94 br_0_94 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c94
*+ bl_0_94 br_0_94 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c94
*+ bl_0_94 br_0_94 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c94
*+ bl_0_94 br_0_94 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c94
*+ bl_0_94 br_0_94 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c94
*+ bl_0_94 br_0_94 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c94
*+ bl_0_94 br_0_94 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c94
*+ bl_0_94 br_0_94 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c94
*+ bl_0_94 br_0_94 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c94
*+ bl_0_94 br_0_94 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c94
*+ bl_0_94 br_0_94 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c94
*+ bl_0_94 br_0_94 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c94
*+ bl_0_94 br_0_94 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c94
*+ bl_0_94 br_0_94 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c94
*+ bl_0_94 br_0_94 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c94
*+ bl_0_94 br_0_94 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c94
*+ bl_0_94 br_0_94 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c94
*+ bl_0_94 br_0_94 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c94
*+ bl_0_94 br_0_94 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c94
*+ bl_0_94 br_0_94 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c94
*+ bl_0_94 br_0_94 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c94
*+ bl_0_94 br_0_94 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c94
*+ bl_0_94 br_0_94 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c94
*+ bl_0_94 br_0_94 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c94
*+ bl_0_94 br_0_94 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c94
*+ bl_0_94 br_0_94 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c94
*+ bl_0_94 br_0_94 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c94
*+ bl_0_94 br_0_94 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c94
*+ bl_0_94 br_0_94 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c94
*+ bl_0_94 br_0_94 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c94
*+ bl_0_94 br_0_94 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c94
*+ bl_0_94 br_0_94 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c94
*+ bl_0_94 br_0_94 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c94
*+ bl_0_94 br_0_94 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c94
*+ bl_0_94 br_0_94 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c94
*+ bl_0_94 br_0_94 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c94
*+ bl_0_94 br_0_94 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c94
*+ bl_0_94 br_0_94 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c94
*+ bl_0_94 br_0_94 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c94
*+ bl_0_94 br_0_94 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c94
*+ bl_0_94 br_0_94 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c94
*+ bl_0_94 br_0_94 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c94
*+ bl_0_94 br_0_94 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c94
*+ bl_0_94 br_0_94 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c94
*+ bl_0_94 br_0_94 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c94
*+ bl_0_94 br_0_94 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c94
*+ bl_0_94 br_0_94 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c94
*+ bl_0_94 br_0_94 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c94
*+ bl_0_94 br_0_94 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c94
*+ bl_0_94 br_0_94 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c94
*+ bl_0_94 br_0_94 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c94
*+ bl_0_94 br_0_94 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c94
*+ bl_0_94 br_0_94 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c94
*+ bl_0_94 br_0_94 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c94
*+ bl_0_94 br_0_94 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c94
*+ bl_0_94 br_0_94 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c94
*+ bl_0_94 br_0_94 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c94
*+ bl_0_94 br_0_94 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c94
*+ bl_0_94 br_0_94 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c94
*+ bl_0_94 br_0_94 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c94
*+ bl_0_94 br_0_94 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c94
*+ bl_0_94 br_0_94 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c94
*+ bl_0_94 br_0_94 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c94
*+ bl_0_94 br_0_94 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c94
*+ bl_0_94 br_0_94 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c94
*+ bl_0_94 br_0_94 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c94
*+ bl_0_94 br_0_94 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c94
*+ bl_0_94 br_0_94 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c94
*+ bl_0_94 br_0_94 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c94
*+ bl_0_94 br_0_94 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c94
*+ bl_0_94 br_0_94 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c94
*+ bl_0_94 br_0_94 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c94
*+ bl_0_94 br_0_94 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c94
*+ bl_0_94 br_0_94 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c94
*+ bl_0_94 br_0_94 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c94
*+ bl_0_94 br_0_94 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c94
*+ bl_0_94 br_0_94 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c94
*+ bl_0_94 br_0_94 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c94
*+ bl_0_94 br_0_94 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c94
*+ bl_0_94 br_0_94 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c94
*+ bl_0_94 br_0_94 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c94
*+ bl_0_94 br_0_94 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c94
*+ bl_0_94 br_0_94 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c94
*+ bl_0_94 br_0_94 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c94
*+ bl_0_94 br_0_94 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c94
*+ bl_0_94 br_0_94 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c94
*+ bl_0_94 br_0_94 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c94
*+ bl_0_94 br_0_94 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c94
*+ bl_0_94 br_0_94 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c94
*+ bl_0_94 br_0_94 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c94
*+ bl_0_94 br_0_94 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c94
*+ bl_0_94 br_0_94 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c94
+ bl_0_94 br_0_94 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c95
+ bl_0_95 br_0_95 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c95
*+ bl_0_95 br_0_95 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c95
*+ bl_0_95 br_0_95 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c95
*+ bl_0_95 br_0_95 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c95
*+ bl_0_95 br_0_95 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c95
*+ bl_0_95 br_0_95 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c95
*+ bl_0_95 br_0_95 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c95
*+ bl_0_95 br_0_95 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c95
*+ bl_0_95 br_0_95 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c95
*+ bl_0_95 br_0_95 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c95
*+ bl_0_95 br_0_95 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c95
*+ bl_0_95 br_0_95 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c95
*+ bl_0_95 br_0_95 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c95
*+ bl_0_95 br_0_95 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c95
*+ bl_0_95 br_0_95 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c95
*+ bl_0_95 br_0_95 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c95
*+ bl_0_95 br_0_95 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c95
*+ bl_0_95 br_0_95 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c95
*+ bl_0_95 br_0_95 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c95
*+ bl_0_95 br_0_95 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c95
*+ bl_0_95 br_0_95 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c95
*+ bl_0_95 br_0_95 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c95
*+ bl_0_95 br_0_95 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c95
*+ bl_0_95 br_0_95 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c95
*+ bl_0_95 br_0_95 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c95
*+ bl_0_95 br_0_95 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c95
*+ bl_0_95 br_0_95 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c95
*+ bl_0_95 br_0_95 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c95
*+ bl_0_95 br_0_95 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c95
*+ bl_0_95 br_0_95 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c95
*+ bl_0_95 br_0_95 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c95
*+ bl_0_95 br_0_95 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c95
*+ bl_0_95 br_0_95 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c95
*+ bl_0_95 br_0_95 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c95
*+ bl_0_95 br_0_95 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c95
*+ bl_0_95 br_0_95 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c95
*+ bl_0_95 br_0_95 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c95
*+ bl_0_95 br_0_95 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c95
*+ bl_0_95 br_0_95 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c95
*+ bl_0_95 br_0_95 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c95
*+ bl_0_95 br_0_95 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c95
*+ bl_0_95 br_0_95 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c95
*+ bl_0_95 br_0_95 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c95
*+ bl_0_95 br_0_95 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c95
*+ bl_0_95 br_0_95 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c95
*+ bl_0_95 br_0_95 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c95
*+ bl_0_95 br_0_95 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c95
*+ bl_0_95 br_0_95 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c95
*+ bl_0_95 br_0_95 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c95
*+ bl_0_95 br_0_95 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c95
*+ bl_0_95 br_0_95 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c95
*+ bl_0_95 br_0_95 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c95
*+ bl_0_95 br_0_95 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c95
*+ bl_0_95 br_0_95 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c95
*+ bl_0_95 br_0_95 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c95
*+ bl_0_95 br_0_95 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c95
*+ bl_0_95 br_0_95 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c95
*+ bl_0_95 br_0_95 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c95
*+ bl_0_95 br_0_95 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c95
*+ bl_0_95 br_0_95 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c95
*+ bl_0_95 br_0_95 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c95
*+ bl_0_95 br_0_95 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c95
*+ bl_0_95 br_0_95 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c95
*+ bl_0_95 br_0_95 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c95
*+ bl_0_95 br_0_95 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c95
*+ bl_0_95 br_0_95 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c95
*+ bl_0_95 br_0_95 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c95
*+ bl_0_95 br_0_95 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c95
*+ bl_0_95 br_0_95 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c95
*+ bl_0_95 br_0_95 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c95
*+ bl_0_95 br_0_95 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c95
*+ bl_0_95 br_0_95 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c95
*+ bl_0_95 br_0_95 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c95
*+ bl_0_95 br_0_95 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c95
*+ bl_0_95 br_0_95 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c95
*+ bl_0_95 br_0_95 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c95
*+ bl_0_95 br_0_95 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c95
*+ bl_0_95 br_0_95 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c95
*+ bl_0_95 br_0_95 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c95
*+ bl_0_95 br_0_95 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c95
*+ bl_0_95 br_0_95 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c95
*+ bl_0_95 br_0_95 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c95
*+ bl_0_95 br_0_95 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c95
*+ bl_0_95 br_0_95 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c95
*+ bl_0_95 br_0_95 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c95
*+ bl_0_95 br_0_95 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c95
*+ bl_0_95 br_0_95 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c95
*+ bl_0_95 br_0_95 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c95
*+ bl_0_95 br_0_95 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c95
*+ bl_0_95 br_0_95 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c95
*+ bl_0_95 br_0_95 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c95
*+ bl_0_95 br_0_95 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c95
*+ bl_0_95 br_0_95 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c95
*+ bl_0_95 br_0_95 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c95
*+ bl_0_95 br_0_95 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c95
*+ bl_0_95 br_0_95 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c95
*+ bl_0_95 br_0_95 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c95
*+ bl_0_95 br_0_95 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c95
*+ bl_0_95 br_0_95 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c95
*+ bl_0_95 br_0_95 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c95
*+ bl_0_95 br_0_95 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c95
*+ bl_0_95 br_0_95 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c95
*+ bl_0_95 br_0_95 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c95
*+ bl_0_95 br_0_95 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c95
*+ bl_0_95 br_0_95 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c95
*+ bl_0_95 br_0_95 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c95
*+ bl_0_95 br_0_95 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c95
*+ bl_0_95 br_0_95 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c95
*+ bl_0_95 br_0_95 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c95
*+ bl_0_95 br_0_95 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c95
*+ bl_0_95 br_0_95 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c95
*+ bl_0_95 br_0_95 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c95
*+ bl_0_95 br_0_95 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c95
*+ bl_0_95 br_0_95 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c95
*+ bl_0_95 br_0_95 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c95
*+ bl_0_95 br_0_95 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c95
*+ bl_0_95 br_0_95 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c95
*+ bl_0_95 br_0_95 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c95
*+ bl_0_95 br_0_95 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c95
*+ bl_0_95 br_0_95 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c95
*+ bl_0_95 br_0_95 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c95
*+ bl_0_95 br_0_95 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c95
*+ bl_0_95 br_0_95 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c95
*+ bl_0_95 br_0_95 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c95
*+ bl_0_95 br_0_95 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c95
*+ bl_0_95 br_0_95 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c95
*+ bl_0_95 br_0_95 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c95
+ bl_0_95 br_0_95 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c96
+ bl_0_96 br_0_96 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c96
*+ bl_0_96 br_0_96 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c96
*+ bl_0_96 br_0_96 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c96
*+ bl_0_96 br_0_96 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c96
*+ bl_0_96 br_0_96 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c96
*+ bl_0_96 br_0_96 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c96
*+ bl_0_96 br_0_96 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c96
*+ bl_0_96 br_0_96 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c96
*+ bl_0_96 br_0_96 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c96
*+ bl_0_96 br_0_96 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c96
*+ bl_0_96 br_0_96 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c96
*+ bl_0_96 br_0_96 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c96
*+ bl_0_96 br_0_96 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c96
*+ bl_0_96 br_0_96 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c96
*+ bl_0_96 br_0_96 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c96
*+ bl_0_96 br_0_96 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c96
*+ bl_0_96 br_0_96 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c96
*+ bl_0_96 br_0_96 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c96
*+ bl_0_96 br_0_96 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c96
*+ bl_0_96 br_0_96 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c96
*+ bl_0_96 br_0_96 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c96
*+ bl_0_96 br_0_96 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c96
*+ bl_0_96 br_0_96 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c96
*+ bl_0_96 br_0_96 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c96
*+ bl_0_96 br_0_96 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c96
*+ bl_0_96 br_0_96 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c96
*+ bl_0_96 br_0_96 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c96
*+ bl_0_96 br_0_96 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c96
*+ bl_0_96 br_0_96 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c96
*+ bl_0_96 br_0_96 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c96
*+ bl_0_96 br_0_96 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c96
*+ bl_0_96 br_0_96 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c96
*+ bl_0_96 br_0_96 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c96
*+ bl_0_96 br_0_96 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c96
*+ bl_0_96 br_0_96 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c96
*+ bl_0_96 br_0_96 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c96
*+ bl_0_96 br_0_96 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c96
*+ bl_0_96 br_0_96 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c96
*+ bl_0_96 br_0_96 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c96
*+ bl_0_96 br_0_96 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c96
*+ bl_0_96 br_0_96 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c96
*+ bl_0_96 br_0_96 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c96
*+ bl_0_96 br_0_96 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c96
*+ bl_0_96 br_0_96 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c96
*+ bl_0_96 br_0_96 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c96
*+ bl_0_96 br_0_96 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c96
*+ bl_0_96 br_0_96 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c96
*+ bl_0_96 br_0_96 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c96
*+ bl_0_96 br_0_96 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c96
*+ bl_0_96 br_0_96 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c96
*+ bl_0_96 br_0_96 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c96
*+ bl_0_96 br_0_96 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c96
*+ bl_0_96 br_0_96 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c96
*+ bl_0_96 br_0_96 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c96
*+ bl_0_96 br_0_96 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c96
*+ bl_0_96 br_0_96 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c96
*+ bl_0_96 br_0_96 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c96
*+ bl_0_96 br_0_96 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c96
*+ bl_0_96 br_0_96 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c96
*+ bl_0_96 br_0_96 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c96
*+ bl_0_96 br_0_96 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c96
*+ bl_0_96 br_0_96 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c96
*+ bl_0_96 br_0_96 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c96
*+ bl_0_96 br_0_96 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c96
*+ bl_0_96 br_0_96 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c96
*+ bl_0_96 br_0_96 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c96
*+ bl_0_96 br_0_96 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c96
*+ bl_0_96 br_0_96 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c96
*+ bl_0_96 br_0_96 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c96
*+ bl_0_96 br_0_96 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c96
*+ bl_0_96 br_0_96 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c96
*+ bl_0_96 br_0_96 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c96
*+ bl_0_96 br_0_96 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c96
*+ bl_0_96 br_0_96 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c96
*+ bl_0_96 br_0_96 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c96
*+ bl_0_96 br_0_96 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c96
*+ bl_0_96 br_0_96 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c96
*+ bl_0_96 br_0_96 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c96
*+ bl_0_96 br_0_96 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c96
*+ bl_0_96 br_0_96 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c96
*+ bl_0_96 br_0_96 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c96
*+ bl_0_96 br_0_96 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c96
*+ bl_0_96 br_0_96 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c96
*+ bl_0_96 br_0_96 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c96
*+ bl_0_96 br_0_96 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c96
*+ bl_0_96 br_0_96 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c96
*+ bl_0_96 br_0_96 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c96
*+ bl_0_96 br_0_96 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c96
*+ bl_0_96 br_0_96 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c96
*+ bl_0_96 br_0_96 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c96
*+ bl_0_96 br_0_96 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c96
*+ bl_0_96 br_0_96 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c96
*+ bl_0_96 br_0_96 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c96
*+ bl_0_96 br_0_96 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c96
*+ bl_0_96 br_0_96 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c96
*+ bl_0_96 br_0_96 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c96
*+ bl_0_96 br_0_96 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c96
*+ bl_0_96 br_0_96 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c96
*+ bl_0_96 br_0_96 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c96
*+ bl_0_96 br_0_96 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c96
*+ bl_0_96 br_0_96 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c96
*+ bl_0_96 br_0_96 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c96
*+ bl_0_96 br_0_96 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c96
*+ bl_0_96 br_0_96 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c96
*+ bl_0_96 br_0_96 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c96
*+ bl_0_96 br_0_96 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c96
*+ bl_0_96 br_0_96 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c96
*+ bl_0_96 br_0_96 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c96
*+ bl_0_96 br_0_96 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c96
*+ bl_0_96 br_0_96 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c96
*+ bl_0_96 br_0_96 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c96
*+ bl_0_96 br_0_96 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c96
*+ bl_0_96 br_0_96 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c96
*+ bl_0_96 br_0_96 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c96
*+ bl_0_96 br_0_96 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c96
*+ bl_0_96 br_0_96 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c96
*+ bl_0_96 br_0_96 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c96
*+ bl_0_96 br_0_96 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c96
*+ bl_0_96 br_0_96 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c96
*+ bl_0_96 br_0_96 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c96
*+ bl_0_96 br_0_96 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c96
*+ bl_0_96 br_0_96 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c96
*+ bl_0_96 br_0_96 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c96
*+ bl_0_96 br_0_96 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c96
*+ bl_0_96 br_0_96 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c96
*+ bl_0_96 br_0_96 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c96
*+ bl_0_96 br_0_96 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c96
+ bl_0_96 br_0_96 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c97
+ bl_0_97 br_0_97 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c97
*+ bl_0_97 br_0_97 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c97
*+ bl_0_97 br_0_97 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c97
*+ bl_0_97 br_0_97 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c97
*+ bl_0_97 br_0_97 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c97
*+ bl_0_97 br_0_97 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c97
*+ bl_0_97 br_0_97 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c97
*+ bl_0_97 br_0_97 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c97
*+ bl_0_97 br_0_97 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c97
*+ bl_0_97 br_0_97 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c97
*+ bl_0_97 br_0_97 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c97
*+ bl_0_97 br_0_97 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c97
*+ bl_0_97 br_0_97 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c97
*+ bl_0_97 br_0_97 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c97
*+ bl_0_97 br_0_97 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c97
*+ bl_0_97 br_0_97 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c97
*+ bl_0_97 br_0_97 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c97
*+ bl_0_97 br_0_97 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c97
*+ bl_0_97 br_0_97 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c97
*+ bl_0_97 br_0_97 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c97
*+ bl_0_97 br_0_97 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c97
*+ bl_0_97 br_0_97 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c97
*+ bl_0_97 br_0_97 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c97
*+ bl_0_97 br_0_97 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c97
*+ bl_0_97 br_0_97 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c97
*+ bl_0_97 br_0_97 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c97
*+ bl_0_97 br_0_97 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c97
*+ bl_0_97 br_0_97 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c97
*+ bl_0_97 br_0_97 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c97
*+ bl_0_97 br_0_97 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c97
*+ bl_0_97 br_0_97 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c97
*+ bl_0_97 br_0_97 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c97
*+ bl_0_97 br_0_97 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c97
*+ bl_0_97 br_0_97 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c97
*+ bl_0_97 br_0_97 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c97
*+ bl_0_97 br_0_97 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c97
*+ bl_0_97 br_0_97 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c97
*+ bl_0_97 br_0_97 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c97
*+ bl_0_97 br_0_97 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c97
*+ bl_0_97 br_0_97 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c97
*+ bl_0_97 br_0_97 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c97
*+ bl_0_97 br_0_97 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c97
*+ bl_0_97 br_0_97 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c97
*+ bl_0_97 br_0_97 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c97
*+ bl_0_97 br_0_97 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c97
*+ bl_0_97 br_0_97 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c97
*+ bl_0_97 br_0_97 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c97
*+ bl_0_97 br_0_97 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c97
*+ bl_0_97 br_0_97 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c97
*+ bl_0_97 br_0_97 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c97
*+ bl_0_97 br_0_97 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c97
*+ bl_0_97 br_0_97 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c97
*+ bl_0_97 br_0_97 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c97
*+ bl_0_97 br_0_97 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c97
*+ bl_0_97 br_0_97 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c97
*+ bl_0_97 br_0_97 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c97
*+ bl_0_97 br_0_97 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c97
*+ bl_0_97 br_0_97 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c97
*+ bl_0_97 br_0_97 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c97
*+ bl_0_97 br_0_97 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c97
*+ bl_0_97 br_0_97 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c97
*+ bl_0_97 br_0_97 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c97
*+ bl_0_97 br_0_97 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c97
*+ bl_0_97 br_0_97 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c97
*+ bl_0_97 br_0_97 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c97
*+ bl_0_97 br_0_97 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c97
*+ bl_0_97 br_0_97 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c97
*+ bl_0_97 br_0_97 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c97
*+ bl_0_97 br_0_97 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c97
*+ bl_0_97 br_0_97 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c97
*+ bl_0_97 br_0_97 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c97
*+ bl_0_97 br_0_97 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c97
*+ bl_0_97 br_0_97 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c97
*+ bl_0_97 br_0_97 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c97
*+ bl_0_97 br_0_97 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c97
*+ bl_0_97 br_0_97 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c97
*+ bl_0_97 br_0_97 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c97
*+ bl_0_97 br_0_97 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c97
*+ bl_0_97 br_0_97 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c97
*+ bl_0_97 br_0_97 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c97
*+ bl_0_97 br_0_97 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c97
*+ bl_0_97 br_0_97 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c97
*+ bl_0_97 br_0_97 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c97
*+ bl_0_97 br_0_97 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c97
*+ bl_0_97 br_0_97 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c97
*+ bl_0_97 br_0_97 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c97
*+ bl_0_97 br_0_97 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c97
*+ bl_0_97 br_0_97 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c97
*+ bl_0_97 br_0_97 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c97
*+ bl_0_97 br_0_97 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c97
*+ bl_0_97 br_0_97 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c97
*+ bl_0_97 br_0_97 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c97
*+ bl_0_97 br_0_97 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c97
*+ bl_0_97 br_0_97 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c97
*+ bl_0_97 br_0_97 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c97
*+ bl_0_97 br_0_97 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c97
*+ bl_0_97 br_0_97 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c97
*+ bl_0_97 br_0_97 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c97
*+ bl_0_97 br_0_97 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c97
*+ bl_0_97 br_0_97 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c97
*+ bl_0_97 br_0_97 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c97
*+ bl_0_97 br_0_97 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c97
*+ bl_0_97 br_0_97 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c97
*+ bl_0_97 br_0_97 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c97
*+ bl_0_97 br_0_97 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c97
*+ bl_0_97 br_0_97 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c97
*+ bl_0_97 br_0_97 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c97
*+ bl_0_97 br_0_97 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c97
*+ bl_0_97 br_0_97 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c97
*+ bl_0_97 br_0_97 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c97
*+ bl_0_97 br_0_97 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c97
*+ bl_0_97 br_0_97 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c97
*+ bl_0_97 br_0_97 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c97
*+ bl_0_97 br_0_97 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c97
*+ bl_0_97 br_0_97 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c97
*+ bl_0_97 br_0_97 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c97
*+ bl_0_97 br_0_97 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c97
*+ bl_0_97 br_0_97 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c97
*+ bl_0_97 br_0_97 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c97
*+ bl_0_97 br_0_97 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c97
*+ bl_0_97 br_0_97 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c97
*+ bl_0_97 br_0_97 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c97
*+ bl_0_97 br_0_97 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c97
*+ bl_0_97 br_0_97 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c97
*+ bl_0_97 br_0_97 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c97
*+ bl_0_97 br_0_97 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c97
*+ bl_0_97 br_0_97 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c97
+ bl_0_97 br_0_97 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c98
+ bl_0_98 br_0_98 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c98
*+ bl_0_98 br_0_98 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c98
*+ bl_0_98 br_0_98 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c98
*+ bl_0_98 br_0_98 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c98
*+ bl_0_98 br_0_98 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c98
*+ bl_0_98 br_0_98 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c98
*+ bl_0_98 br_0_98 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c98
*+ bl_0_98 br_0_98 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c98
*+ bl_0_98 br_0_98 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c98
*+ bl_0_98 br_0_98 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c98
*+ bl_0_98 br_0_98 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c98
*+ bl_0_98 br_0_98 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c98
*+ bl_0_98 br_0_98 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c98
*+ bl_0_98 br_0_98 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c98
*+ bl_0_98 br_0_98 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c98
*+ bl_0_98 br_0_98 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c98
*+ bl_0_98 br_0_98 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c98
*+ bl_0_98 br_0_98 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c98
*+ bl_0_98 br_0_98 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c98
*+ bl_0_98 br_0_98 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c98
*+ bl_0_98 br_0_98 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c98
*+ bl_0_98 br_0_98 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c98
*+ bl_0_98 br_0_98 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c98
*+ bl_0_98 br_0_98 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c98
*+ bl_0_98 br_0_98 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c98
*+ bl_0_98 br_0_98 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c98
*+ bl_0_98 br_0_98 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c98
*+ bl_0_98 br_0_98 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c98
*+ bl_0_98 br_0_98 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c98
*+ bl_0_98 br_0_98 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c98
*+ bl_0_98 br_0_98 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c98
*+ bl_0_98 br_0_98 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c98
*+ bl_0_98 br_0_98 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c98
*+ bl_0_98 br_0_98 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c98
*+ bl_0_98 br_0_98 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c98
*+ bl_0_98 br_0_98 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c98
*+ bl_0_98 br_0_98 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c98
*+ bl_0_98 br_0_98 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c98
*+ bl_0_98 br_0_98 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c98
*+ bl_0_98 br_0_98 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c98
*+ bl_0_98 br_0_98 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c98
*+ bl_0_98 br_0_98 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c98
*+ bl_0_98 br_0_98 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c98
*+ bl_0_98 br_0_98 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c98
*+ bl_0_98 br_0_98 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c98
*+ bl_0_98 br_0_98 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c98
*+ bl_0_98 br_0_98 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c98
*+ bl_0_98 br_0_98 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c98
*+ bl_0_98 br_0_98 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c98
*+ bl_0_98 br_0_98 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c98
*+ bl_0_98 br_0_98 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c98
*+ bl_0_98 br_0_98 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c98
*+ bl_0_98 br_0_98 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c98
*+ bl_0_98 br_0_98 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c98
*+ bl_0_98 br_0_98 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c98
*+ bl_0_98 br_0_98 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c98
*+ bl_0_98 br_0_98 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c98
*+ bl_0_98 br_0_98 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c98
*+ bl_0_98 br_0_98 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c98
*+ bl_0_98 br_0_98 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c98
*+ bl_0_98 br_0_98 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c98
*+ bl_0_98 br_0_98 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c98
*+ bl_0_98 br_0_98 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c98
*+ bl_0_98 br_0_98 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c98
*+ bl_0_98 br_0_98 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c98
*+ bl_0_98 br_0_98 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c98
*+ bl_0_98 br_0_98 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c98
*+ bl_0_98 br_0_98 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c98
*+ bl_0_98 br_0_98 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c98
*+ bl_0_98 br_0_98 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c98
*+ bl_0_98 br_0_98 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c98
*+ bl_0_98 br_0_98 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c98
*+ bl_0_98 br_0_98 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c98
*+ bl_0_98 br_0_98 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c98
*+ bl_0_98 br_0_98 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c98
*+ bl_0_98 br_0_98 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c98
*+ bl_0_98 br_0_98 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c98
*+ bl_0_98 br_0_98 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c98
*+ bl_0_98 br_0_98 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c98
*+ bl_0_98 br_0_98 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c98
*+ bl_0_98 br_0_98 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c98
*+ bl_0_98 br_0_98 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c98
*+ bl_0_98 br_0_98 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c98
*+ bl_0_98 br_0_98 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c98
*+ bl_0_98 br_0_98 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c98
*+ bl_0_98 br_0_98 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c98
*+ bl_0_98 br_0_98 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c98
*+ bl_0_98 br_0_98 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c98
*+ bl_0_98 br_0_98 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c98
*+ bl_0_98 br_0_98 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c98
*+ bl_0_98 br_0_98 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c98
*+ bl_0_98 br_0_98 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c98
*+ bl_0_98 br_0_98 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c98
*+ bl_0_98 br_0_98 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c98
*+ bl_0_98 br_0_98 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c98
*+ bl_0_98 br_0_98 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c98
*+ bl_0_98 br_0_98 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c98
*+ bl_0_98 br_0_98 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c98
*+ bl_0_98 br_0_98 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c98
*+ bl_0_98 br_0_98 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c98
*+ bl_0_98 br_0_98 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c98
*+ bl_0_98 br_0_98 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c98
*+ bl_0_98 br_0_98 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c98
*+ bl_0_98 br_0_98 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c98
*+ bl_0_98 br_0_98 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c98
*+ bl_0_98 br_0_98 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c98
*+ bl_0_98 br_0_98 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c98
*+ bl_0_98 br_0_98 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c98
*+ bl_0_98 br_0_98 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c98
*+ bl_0_98 br_0_98 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c98
*+ bl_0_98 br_0_98 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c98
*+ bl_0_98 br_0_98 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c98
*+ bl_0_98 br_0_98 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c98
*+ bl_0_98 br_0_98 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c98
*+ bl_0_98 br_0_98 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c98
*+ bl_0_98 br_0_98 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c98
*+ bl_0_98 br_0_98 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c98
*+ bl_0_98 br_0_98 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c98
*+ bl_0_98 br_0_98 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c98
*+ bl_0_98 br_0_98 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c98
*+ bl_0_98 br_0_98 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c98
*+ bl_0_98 br_0_98 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c98
*+ bl_0_98 br_0_98 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c98
*+ bl_0_98 br_0_98 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c98
*+ bl_0_98 br_0_98 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c98
*+ bl_0_98 br_0_98 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c98
*+ bl_0_98 br_0_98 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c98
+ bl_0_98 br_0_98 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c99
+ bl_0_99 br_0_99 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c99
*+ bl_0_99 br_0_99 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c99
*+ bl_0_99 br_0_99 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c99
*+ bl_0_99 br_0_99 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c99
*+ bl_0_99 br_0_99 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c99
*+ bl_0_99 br_0_99 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c99
*+ bl_0_99 br_0_99 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c99
*+ bl_0_99 br_0_99 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c99
*+ bl_0_99 br_0_99 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c99
*+ bl_0_99 br_0_99 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c99
*+ bl_0_99 br_0_99 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c99
*+ bl_0_99 br_0_99 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c99
*+ bl_0_99 br_0_99 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c99
*+ bl_0_99 br_0_99 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c99
*+ bl_0_99 br_0_99 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c99
*+ bl_0_99 br_0_99 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c99
*+ bl_0_99 br_0_99 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c99
*+ bl_0_99 br_0_99 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c99
*+ bl_0_99 br_0_99 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c99
*+ bl_0_99 br_0_99 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c99
*+ bl_0_99 br_0_99 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c99
*+ bl_0_99 br_0_99 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c99
*+ bl_0_99 br_0_99 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c99
*+ bl_0_99 br_0_99 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c99
*+ bl_0_99 br_0_99 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c99
*+ bl_0_99 br_0_99 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c99
*+ bl_0_99 br_0_99 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c99
*+ bl_0_99 br_0_99 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c99
*+ bl_0_99 br_0_99 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c99
*+ bl_0_99 br_0_99 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c99
*+ bl_0_99 br_0_99 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c99
*+ bl_0_99 br_0_99 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c99
*+ bl_0_99 br_0_99 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c99
*+ bl_0_99 br_0_99 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c99
*+ bl_0_99 br_0_99 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c99
*+ bl_0_99 br_0_99 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c99
*+ bl_0_99 br_0_99 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c99
*+ bl_0_99 br_0_99 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c99
*+ bl_0_99 br_0_99 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c99
*+ bl_0_99 br_0_99 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c99
*+ bl_0_99 br_0_99 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c99
*+ bl_0_99 br_0_99 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c99
*+ bl_0_99 br_0_99 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c99
*+ bl_0_99 br_0_99 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c99
*+ bl_0_99 br_0_99 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c99
*+ bl_0_99 br_0_99 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c99
*+ bl_0_99 br_0_99 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c99
*+ bl_0_99 br_0_99 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c99
*+ bl_0_99 br_0_99 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c99
*+ bl_0_99 br_0_99 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c99
*+ bl_0_99 br_0_99 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c99
*+ bl_0_99 br_0_99 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c99
*+ bl_0_99 br_0_99 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c99
*+ bl_0_99 br_0_99 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c99
*+ bl_0_99 br_0_99 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c99
*+ bl_0_99 br_0_99 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c99
*+ bl_0_99 br_0_99 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c99
*+ bl_0_99 br_0_99 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c99
*+ bl_0_99 br_0_99 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c99
*+ bl_0_99 br_0_99 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c99
*+ bl_0_99 br_0_99 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c99
*+ bl_0_99 br_0_99 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c99
*+ bl_0_99 br_0_99 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c99
*+ bl_0_99 br_0_99 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c99
*+ bl_0_99 br_0_99 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c99
*+ bl_0_99 br_0_99 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c99
*+ bl_0_99 br_0_99 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c99
*+ bl_0_99 br_0_99 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c99
*+ bl_0_99 br_0_99 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c99
*+ bl_0_99 br_0_99 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c99
*+ bl_0_99 br_0_99 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c99
*+ bl_0_99 br_0_99 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c99
*+ bl_0_99 br_0_99 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c99
*+ bl_0_99 br_0_99 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c99
*+ bl_0_99 br_0_99 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c99
*+ bl_0_99 br_0_99 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c99
*+ bl_0_99 br_0_99 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c99
*+ bl_0_99 br_0_99 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c99
*+ bl_0_99 br_0_99 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c99
*+ bl_0_99 br_0_99 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c99
*+ bl_0_99 br_0_99 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c99
*+ bl_0_99 br_0_99 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c99
*+ bl_0_99 br_0_99 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c99
*+ bl_0_99 br_0_99 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c99
*+ bl_0_99 br_0_99 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c99
*+ bl_0_99 br_0_99 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c99
*+ bl_0_99 br_0_99 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c99
*+ bl_0_99 br_0_99 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c99
*+ bl_0_99 br_0_99 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c99
*+ bl_0_99 br_0_99 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c99
*+ bl_0_99 br_0_99 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c99
*+ bl_0_99 br_0_99 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c99
*+ bl_0_99 br_0_99 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c99
*+ bl_0_99 br_0_99 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c99
*+ bl_0_99 br_0_99 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c99
*+ bl_0_99 br_0_99 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c99
*+ bl_0_99 br_0_99 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c99
*+ bl_0_99 br_0_99 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c99
*+ bl_0_99 br_0_99 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c99
*+ bl_0_99 br_0_99 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c99
*+ bl_0_99 br_0_99 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c99
*+ bl_0_99 br_0_99 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c99
*+ bl_0_99 br_0_99 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c99
*+ bl_0_99 br_0_99 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c99
*+ bl_0_99 br_0_99 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c99
*+ bl_0_99 br_0_99 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c99
*+ bl_0_99 br_0_99 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c99
*+ bl_0_99 br_0_99 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c99
*+ bl_0_99 br_0_99 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c99
*+ bl_0_99 br_0_99 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c99
*+ bl_0_99 br_0_99 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c99
*+ bl_0_99 br_0_99 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c99
*+ bl_0_99 br_0_99 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c99
*+ bl_0_99 br_0_99 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c99
*+ bl_0_99 br_0_99 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c99
*+ bl_0_99 br_0_99 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c99
*+ bl_0_99 br_0_99 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c99
*+ bl_0_99 br_0_99 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c99
*+ bl_0_99 br_0_99 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c99
*+ bl_0_99 br_0_99 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c99
*+ bl_0_99 br_0_99 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c99
*+ bl_0_99 br_0_99 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c99
*+ bl_0_99 br_0_99 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c99
*+ bl_0_99 br_0_99 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c99
*+ bl_0_99 br_0_99 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c99
*+ bl_0_99 br_0_99 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c99
*+ bl_0_99 br_0_99 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c99
+ bl_0_99 br_0_99 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c100
+ bl_0_100 br_0_100 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c100
*+ bl_0_100 br_0_100 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c100
*+ bl_0_100 br_0_100 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c100
*+ bl_0_100 br_0_100 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c100
*+ bl_0_100 br_0_100 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c100
*+ bl_0_100 br_0_100 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c100
*+ bl_0_100 br_0_100 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c100
*+ bl_0_100 br_0_100 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c100
*+ bl_0_100 br_0_100 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c100
*+ bl_0_100 br_0_100 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c100
*+ bl_0_100 br_0_100 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c100
*+ bl_0_100 br_0_100 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c100
*+ bl_0_100 br_0_100 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c100
*+ bl_0_100 br_0_100 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c100
*+ bl_0_100 br_0_100 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c100
*+ bl_0_100 br_0_100 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c100
*+ bl_0_100 br_0_100 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c100
*+ bl_0_100 br_0_100 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c100
*+ bl_0_100 br_0_100 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c100
*+ bl_0_100 br_0_100 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c100
*+ bl_0_100 br_0_100 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c100
*+ bl_0_100 br_0_100 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c100
*+ bl_0_100 br_0_100 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c100
*+ bl_0_100 br_0_100 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c100
*+ bl_0_100 br_0_100 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c100
*+ bl_0_100 br_0_100 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c100
*+ bl_0_100 br_0_100 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c100
*+ bl_0_100 br_0_100 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c100
*+ bl_0_100 br_0_100 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c100
*+ bl_0_100 br_0_100 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c100
*+ bl_0_100 br_0_100 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c100
*+ bl_0_100 br_0_100 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c100
*+ bl_0_100 br_0_100 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c100
*+ bl_0_100 br_0_100 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c100
*+ bl_0_100 br_0_100 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c100
*+ bl_0_100 br_0_100 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c100
*+ bl_0_100 br_0_100 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c100
*+ bl_0_100 br_0_100 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c100
*+ bl_0_100 br_0_100 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c100
*+ bl_0_100 br_0_100 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c100
*+ bl_0_100 br_0_100 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c100
*+ bl_0_100 br_0_100 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c100
*+ bl_0_100 br_0_100 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c100
*+ bl_0_100 br_0_100 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c100
*+ bl_0_100 br_0_100 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c100
*+ bl_0_100 br_0_100 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c100
*+ bl_0_100 br_0_100 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c100
*+ bl_0_100 br_0_100 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c100
*+ bl_0_100 br_0_100 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c100
*+ bl_0_100 br_0_100 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c100
*+ bl_0_100 br_0_100 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c100
*+ bl_0_100 br_0_100 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c100
*+ bl_0_100 br_0_100 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c100
*+ bl_0_100 br_0_100 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c100
*+ bl_0_100 br_0_100 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c100
*+ bl_0_100 br_0_100 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c100
*+ bl_0_100 br_0_100 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c100
*+ bl_0_100 br_0_100 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c100
*+ bl_0_100 br_0_100 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c100
*+ bl_0_100 br_0_100 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c100
*+ bl_0_100 br_0_100 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c100
*+ bl_0_100 br_0_100 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c100
*+ bl_0_100 br_0_100 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c100
*+ bl_0_100 br_0_100 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c100
*+ bl_0_100 br_0_100 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c100
*+ bl_0_100 br_0_100 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c100
*+ bl_0_100 br_0_100 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c100
*+ bl_0_100 br_0_100 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c100
*+ bl_0_100 br_0_100 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c100
*+ bl_0_100 br_0_100 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c100
*+ bl_0_100 br_0_100 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c100
*+ bl_0_100 br_0_100 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c100
*+ bl_0_100 br_0_100 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c100
*+ bl_0_100 br_0_100 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c100
*+ bl_0_100 br_0_100 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c100
*+ bl_0_100 br_0_100 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c100
*+ bl_0_100 br_0_100 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c100
*+ bl_0_100 br_0_100 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c100
*+ bl_0_100 br_0_100 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c100
*+ bl_0_100 br_0_100 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c100
*+ bl_0_100 br_0_100 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c100
*+ bl_0_100 br_0_100 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c100
*+ bl_0_100 br_0_100 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c100
*+ bl_0_100 br_0_100 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c100
*+ bl_0_100 br_0_100 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c100
*+ bl_0_100 br_0_100 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c100
*+ bl_0_100 br_0_100 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c100
*+ bl_0_100 br_0_100 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c100
*+ bl_0_100 br_0_100 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c100
*+ bl_0_100 br_0_100 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c100
*+ bl_0_100 br_0_100 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c100
*+ bl_0_100 br_0_100 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c100
*+ bl_0_100 br_0_100 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c100
*+ bl_0_100 br_0_100 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c100
*+ bl_0_100 br_0_100 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c100
*+ bl_0_100 br_0_100 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c100
*+ bl_0_100 br_0_100 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c100
*+ bl_0_100 br_0_100 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c100
*+ bl_0_100 br_0_100 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c100
*+ bl_0_100 br_0_100 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c100
*+ bl_0_100 br_0_100 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c100
*+ bl_0_100 br_0_100 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c100
*+ bl_0_100 br_0_100 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c100
*+ bl_0_100 br_0_100 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c100
*+ bl_0_100 br_0_100 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c100
*+ bl_0_100 br_0_100 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c100
*+ bl_0_100 br_0_100 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c100
*+ bl_0_100 br_0_100 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c100
*+ bl_0_100 br_0_100 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c100
*+ bl_0_100 br_0_100 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c100
*+ bl_0_100 br_0_100 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c100
*+ bl_0_100 br_0_100 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c100
*+ bl_0_100 br_0_100 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c100
*+ bl_0_100 br_0_100 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c100
*+ bl_0_100 br_0_100 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c100
*+ bl_0_100 br_0_100 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c100
*+ bl_0_100 br_0_100 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c100
*+ bl_0_100 br_0_100 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c100
*+ bl_0_100 br_0_100 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c100
*+ bl_0_100 br_0_100 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c100
*+ bl_0_100 br_0_100 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c100
*+ bl_0_100 br_0_100 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c100
*+ bl_0_100 br_0_100 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c100
*+ bl_0_100 br_0_100 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c100
*+ bl_0_100 br_0_100 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c100
*+ bl_0_100 br_0_100 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c100
*+ bl_0_100 br_0_100 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c100
+ bl_0_100 br_0_100 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c101
+ bl_0_101 br_0_101 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c101
*+ bl_0_101 br_0_101 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c101
*+ bl_0_101 br_0_101 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c101
*+ bl_0_101 br_0_101 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c101
*+ bl_0_101 br_0_101 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c101
*+ bl_0_101 br_0_101 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c101
*+ bl_0_101 br_0_101 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c101
*+ bl_0_101 br_0_101 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c101
*+ bl_0_101 br_0_101 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c101
*+ bl_0_101 br_0_101 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c101
*+ bl_0_101 br_0_101 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c101
*+ bl_0_101 br_0_101 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c101
*+ bl_0_101 br_0_101 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c101
*+ bl_0_101 br_0_101 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c101
*+ bl_0_101 br_0_101 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c101
*+ bl_0_101 br_0_101 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c101
*+ bl_0_101 br_0_101 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c101
*+ bl_0_101 br_0_101 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c101
*+ bl_0_101 br_0_101 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c101
*+ bl_0_101 br_0_101 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c101
*+ bl_0_101 br_0_101 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c101
*+ bl_0_101 br_0_101 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c101
*+ bl_0_101 br_0_101 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c101
*+ bl_0_101 br_0_101 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c101
*+ bl_0_101 br_0_101 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c101
*+ bl_0_101 br_0_101 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c101
*+ bl_0_101 br_0_101 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c101
*+ bl_0_101 br_0_101 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c101
*+ bl_0_101 br_0_101 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c101
*+ bl_0_101 br_0_101 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c101
*+ bl_0_101 br_0_101 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c101
*+ bl_0_101 br_0_101 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c101
*+ bl_0_101 br_0_101 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c101
*+ bl_0_101 br_0_101 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c101
*+ bl_0_101 br_0_101 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c101
*+ bl_0_101 br_0_101 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c101
*+ bl_0_101 br_0_101 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c101
*+ bl_0_101 br_0_101 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c101
*+ bl_0_101 br_0_101 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c101
*+ bl_0_101 br_0_101 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c101
*+ bl_0_101 br_0_101 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c101
*+ bl_0_101 br_0_101 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c101
*+ bl_0_101 br_0_101 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c101
*+ bl_0_101 br_0_101 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c101
*+ bl_0_101 br_0_101 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c101
*+ bl_0_101 br_0_101 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c101
*+ bl_0_101 br_0_101 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c101
*+ bl_0_101 br_0_101 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c101
*+ bl_0_101 br_0_101 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c101
*+ bl_0_101 br_0_101 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c101
*+ bl_0_101 br_0_101 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c101
*+ bl_0_101 br_0_101 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c101
*+ bl_0_101 br_0_101 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c101
*+ bl_0_101 br_0_101 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c101
*+ bl_0_101 br_0_101 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c101
*+ bl_0_101 br_0_101 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c101
*+ bl_0_101 br_0_101 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c101
*+ bl_0_101 br_0_101 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c101
*+ bl_0_101 br_0_101 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c101
*+ bl_0_101 br_0_101 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c101
*+ bl_0_101 br_0_101 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c101
*+ bl_0_101 br_0_101 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c101
*+ bl_0_101 br_0_101 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c101
*+ bl_0_101 br_0_101 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c101
*+ bl_0_101 br_0_101 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c101
*+ bl_0_101 br_0_101 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c101
*+ bl_0_101 br_0_101 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c101
*+ bl_0_101 br_0_101 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c101
*+ bl_0_101 br_0_101 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c101
*+ bl_0_101 br_0_101 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c101
*+ bl_0_101 br_0_101 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c101
*+ bl_0_101 br_0_101 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c101
*+ bl_0_101 br_0_101 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c101
*+ bl_0_101 br_0_101 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c101
*+ bl_0_101 br_0_101 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c101
*+ bl_0_101 br_0_101 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c101
*+ bl_0_101 br_0_101 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c101
*+ bl_0_101 br_0_101 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c101
*+ bl_0_101 br_0_101 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c101
*+ bl_0_101 br_0_101 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c101
*+ bl_0_101 br_0_101 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c101
*+ bl_0_101 br_0_101 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c101
*+ bl_0_101 br_0_101 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c101
*+ bl_0_101 br_0_101 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c101
*+ bl_0_101 br_0_101 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c101
*+ bl_0_101 br_0_101 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c101
*+ bl_0_101 br_0_101 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c101
*+ bl_0_101 br_0_101 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c101
*+ bl_0_101 br_0_101 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c101
*+ bl_0_101 br_0_101 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c101
*+ bl_0_101 br_0_101 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c101
*+ bl_0_101 br_0_101 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c101
*+ bl_0_101 br_0_101 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c101
*+ bl_0_101 br_0_101 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c101
*+ bl_0_101 br_0_101 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c101
*+ bl_0_101 br_0_101 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c101
*+ bl_0_101 br_0_101 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c101
*+ bl_0_101 br_0_101 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c101
*+ bl_0_101 br_0_101 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c101
*+ bl_0_101 br_0_101 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c101
*+ bl_0_101 br_0_101 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c101
*+ bl_0_101 br_0_101 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c101
*+ bl_0_101 br_0_101 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c101
*+ bl_0_101 br_0_101 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c101
*+ bl_0_101 br_0_101 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c101
*+ bl_0_101 br_0_101 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c101
*+ bl_0_101 br_0_101 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c101
*+ bl_0_101 br_0_101 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c101
*+ bl_0_101 br_0_101 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c101
*+ bl_0_101 br_0_101 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c101
*+ bl_0_101 br_0_101 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c101
*+ bl_0_101 br_0_101 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c101
*+ bl_0_101 br_0_101 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c101
*+ bl_0_101 br_0_101 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c101
*+ bl_0_101 br_0_101 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c101
*+ bl_0_101 br_0_101 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c101
*+ bl_0_101 br_0_101 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c101
*+ bl_0_101 br_0_101 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c101
*+ bl_0_101 br_0_101 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c101
*+ bl_0_101 br_0_101 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c101
*+ bl_0_101 br_0_101 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c101
*+ bl_0_101 br_0_101 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c101
*+ bl_0_101 br_0_101 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c101
*+ bl_0_101 br_0_101 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c101
*+ bl_0_101 br_0_101 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c101
*+ bl_0_101 br_0_101 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c101
*+ bl_0_101 br_0_101 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c101
+ bl_0_101 br_0_101 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c102
+ bl_0_102 br_0_102 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c102
*+ bl_0_102 br_0_102 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c102
*+ bl_0_102 br_0_102 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c102
*+ bl_0_102 br_0_102 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c102
*+ bl_0_102 br_0_102 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c102
*+ bl_0_102 br_0_102 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c102
*+ bl_0_102 br_0_102 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c102
*+ bl_0_102 br_0_102 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c102
*+ bl_0_102 br_0_102 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c102
*+ bl_0_102 br_0_102 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c102
*+ bl_0_102 br_0_102 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c102
*+ bl_0_102 br_0_102 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c102
*+ bl_0_102 br_0_102 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c102
*+ bl_0_102 br_0_102 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c102
*+ bl_0_102 br_0_102 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c102
*+ bl_0_102 br_0_102 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c102
*+ bl_0_102 br_0_102 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c102
*+ bl_0_102 br_0_102 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c102
*+ bl_0_102 br_0_102 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c102
*+ bl_0_102 br_0_102 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c102
*+ bl_0_102 br_0_102 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c102
*+ bl_0_102 br_0_102 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c102
*+ bl_0_102 br_0_102 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c102
*+ bl_0_102 br_0_102 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c102
*+ bl_0_102 br_0_102 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c102
*+ bl_0_102 br_0_102 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c102
*+ bl_0_102 br_0_102 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c102
*+ bl_0_102 br_0_102 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c102
*+ bl_0_102 br_0_102 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c102
*+ bl_0_102 br_0_102 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c102
*+ bl_0_102 br_0_102 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c102
*+ bl_0_102 br_0_102 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c102
*+ bl_0_102 br_0_102 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c102
*+ bl_0_102 br_0_102 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c102
*+ bl_0_102 br_0_102 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c102
*+ bl_0_102 br_0_102 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c102
*+ bl_0_102 br_0_102 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c102
*+ bl_0_102 br_0_102 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c102
*+ bl_0_102 br_0_102 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c102
*+ bl_0_102 br_0_102 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c102
*+ bl_0_102 br_0_102 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c102
*+ bl_0_102 br_0_102 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c102
*+ bl_0_102 br_0_102 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c102
*+ bl_0_102 br_0_102 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c102
*+ bl_0_102 br_0_102 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c102
*+ bl_0_102 br_0_102 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c102
*+ bl_0_102 br_0_102 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c102
*+ bl_0_102 br_0_102 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c102
*+ bl_0_102 br_0_102 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c102
*+ bl_0_102 br_0_102 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c102
*+ bl_0_102 br_0_102 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c102
*+ bl_0_102 br_0_102 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c102
*+ bl_0_102 br_0_102 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c102
*+ bl_0_102 br_0_102 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c102
*+ bl_0_102 br_0_102 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c102
*+ bl_0_102 br_0_102 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c102
*+ bl_0_102 br_0_102 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c102
*+ bl_0_102 br_0_102 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c102
*+ bl_0_102 br_0_102 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c102
*+ bl_0_102 br_0_102 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c102
*+ bl_0_102 br_0_102 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c102
*+ bl_0_102 br_0_102 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c102
*+ bl_0_102 br_0_102 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c102
*+ bl_0_102 br_0_102 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c102
*+ bl_0_102 br_0_102 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c102
*+ bl_0_102 br_0_102 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c102
*+ bl_0_102 br_0_102 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c102
*+ bl_0_102 br_0_102 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c102
*+ bl_0_102 br_0_102 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c102
*+ bl_0_102 br_0_102 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c102
*+ bl_0_102 br_0_102 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c102
*+ bl_0_102 br_0_102 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c102
*+ bl_0_102 br_0_102 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c102
*+ bl_0_102 br_0_102 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c102
*+ bl_0_102 br_0_102 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c102
*+ bl_0_102 br_0_102 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c102
*+ bl_0_102 br_0_102 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c102
*+ bl_0_102 br_0_102 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c102
*+ bl_0_102 br_0_102 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c102
*+ bl_0_102 br_0_102 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c102
*+ bl_0_102 br_0_102 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c102
*+ bl_0_102 br_0_102 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c102
*+ bl_0_102 br_0_102 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c102
*+ bl_0_102 br_0_102 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c102
*+ bl_0_102 br_0_102 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c102
*+ bl_0_102 br_0_102 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c102
*+ bl_0_102 br_0_102 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c102
*+ bl_0_102 br_0_102 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c102
*+ bl_0_102 br_0_102 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c102
*+ bl_0_102 br_0_102 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c102
*+ bl_0_102 br_0_102 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c102
*+ bl_0_102 br_0_102 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c102
*+ bl_0_102 br_0_102 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c102
*+ bl_0_102 br_0_102 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c102
*+ bl_0_102 br_0_102 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c102
*+ bl_0_102 br_0_102 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c102
*+ bl_0_102 br_0_102 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c102
*+ bl_0_102 br_0_102 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c102
*+ bl_0_102 br_0_102 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c102
*+ bl_0_102 br_0_102 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c102
*+ bl_0_102 br_0_102 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c102
*+ bl_0_102 br_0_102 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c102
*+ bl_0_102 br_0_102 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c102
*+ bl_0_102 br_0_102 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c102
*+ bl_0_102 br_0_102 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c102
*+ bl_0_102 br_0_102 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c102
*+ bl_0_102 br_0_102 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c102
*+ bl_0_102 br_0_102 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c102
*+ bl_0_102 br_0_102 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c102
*+ bl_0_102 br_0_102 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c102
*+ bl_0_102 br_0_102 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c102
*+ bl_0_102 br_0_102 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c102
*+ bl_0_102 br_0_102 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c102
*+ bl_0_102 br_0_102 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c102
*+ bl_0_102 br_0_102 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c102
*+ bl_0_102 br_0_102 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c102
*+ bl_0_102 br_0_102 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c102
*+ bl_0_102 br_0_102 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c102
*+ bl_0_102 br_0_102 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c102
*+ bl_0_102 br_0_102 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c102
*+ bl_0_102 br_0_102 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c102
*+ bl_0_102 br_0_102 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c102
*+ bl_0_102 br_0_102 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c102
*+ bl_0_102 br_0_102 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c102
*+ bl_0_102 br_0_102 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c102
*+ bl_0_102 br_0_102 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c102
*+ bl_0_102 br_0_102 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c102
+ bl_0_102 br_0_102 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c103
+ bl_0_103 br_0_103 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c103
*+ bl_0_103 br_0_103 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c103
*+ bl_0_103 br_0_103 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c103
*+ bl_0_103 br_0_103 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c103
*+ bl_0_103 br_0_103 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c103
*+ bl_0_103 br_0_103 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c103
*+ bl_0_103 br_0_103 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c103
*+ bl_0_103 br_0_103 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c103
*+ bl_0_103 br_0_103 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c103
*+ bl_0_103 br_0_103 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c103
*+ bl_0_103 br_0_103 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c103
*+ bl_0_103 br_0_103 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c103
*+ bl_0_103 br_0_103 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c103
*+ bl_0_103 br_0_103 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c103
*+ bl_0_103 br_0_103 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c103
*+ bl_0_103 br_0_103 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c103
*+ bl_0_103 br_0_103 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c103
*+ bl_0_103 br_0_103 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c103
*+ bl_0_103 br_0_103 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c103
*+ bl_0_103 br_0_103 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c103
*+ bl_0_103 br_0_103 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c103
*+ bl_0_103 br_0_103 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c103
*+ bl_0_103 br_0_103 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c103
*+ bl_0_103 br_0_103 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c103
*+ bl_0_103 br_0_103 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c103
*+ bl_0_103 br_0_103 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c103
*+ bl_0_103 br_0_103 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c103
*+ bl_0_103 br_0_103 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c103
*+ bl_0_103 br_0_103 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c103
*+ bl_0_103 br_0_103 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c103
*+ bl_0_103 br_0_103 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c103
*+ bl_0_103 br_0_103 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c103
*+ bl_0_103 br_0_103 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c103
*+ bl_0_103 br_0_103 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c103
*+ bl_0_103 br_0_103 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c103
*+ bl_0_103 br_0_103 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c103
*+ bl_0_103 br_0_103 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c103
*+ bl_0_103 br_0_103 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c103
*+ bl_0_103 br_0_103 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c103
*+ bl_0_103 br_0_103 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c103
*+ bl_0_103 br_0_103 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c103
*+ bl_0_103 br_0_103 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c103
*+ bl_0_103 br_0_103 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c103
*+ bl_0_103 br_0_103 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c103
*+ bl_0_103 br_0_103 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c103
*+ bl_0_103 br_0_103 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c103
*+ bl_0_103 br_0_103 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c103
*+ bl_0_103 br_0_103 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c103
*+ bl_0_103 br_0_103 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c103
*+ bl_0_103 br_0_103 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c103
*+ bl_0_103 br_0_103 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c103
*+ bl_0_103 br_0_103 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c103
*+ bl_0_103 br_0_103 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c103
*+ bl_0_103 br_0_103 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c103
*+ bl_0_103 br_0_103 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c103
*+ bl_0_103 br_0_103 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c103
*+ bl_0_103 br_0_103 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c103
*+ bl_0_103 br_0_103 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c103
*+ bl_0_103 br_0_103 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c103
*+ bl_0_103 br_0_103 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c103
*+ bl_0_103 br_0_103 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c103
*+ bl_0_103 br_0_103 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c103
*+ bl_0_103 br_0_103 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c103
*+ bl_0_103 br_0_103 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c103
*+ bl_0_103 br_0_103 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c103
*+ bl_0_103 br_0_103 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c103
*+ bl_0_103 br_0_103 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c103
*+ bl_0_103 br_0_103 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c103
*+ bl_0_103 br_0_103 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c103
*+ bl_0_103 br_0_103 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c103
*+ bl_0_103 br_0_103 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c103
*+ bl_0_103 br_0_103 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c103
*+ bl_0_103 br_0_103 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c103
*+ bl_0_103 br_0_103 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c103
*+ bl_0_103 br_0_103 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c103
*+ bl_0_103 br_0_103 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c103
*+ bl_0_103 br_0_103 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c103
*+ bl_0_103 br_0_103 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c103
*+ bl_0_103 br_0_103 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c103
*+ bl_0_103 br_0_103 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c103
*+ bl_0_103 br_0_103 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c103
*+ bl_0_103 br_0_103 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c103
*+ bl_0_103 br_0_103 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c103
*+ bl_0_103 br_0_103 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c103
*+ bl_0_103 br_0_103 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c103
*+ bl_0_103 br_0_103 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c103
*+ bl_0_103 br_0_103 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c103
*+ bl_0_103 br_0_103 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c103
*+ bl_0_103 br_0_103 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c103
*+ bl_0_103 br_0_103 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c103
*+ bl_0_103 br_0_103 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c103
*+ bl_0_103 br_0_103 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c103
*+ bl_0_103 br_0_103 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c103
*+ bl_0_103 br_0_103 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c103
*+ bl_0_103 br_0_103 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c103
*+ bl_0_103 br_0_103 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c103
*+ bl_0_103 br_0_103 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c103
*+ bl_0_103 br_0_103 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c103
*+ bl_0_103 br_0_103 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c103
*+ bl_0_103 br_0_103 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c103
*+ bl_0_103 br_0_103 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c103
*+ bl_0_103 br_0_103 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c103
*+ bl_0_103 br_0_103 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c103
*+ bl_0_103 br_0_103 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c103
*+ bl_0_103 br_0_103 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c103
*+ bl_0_103 br_0_103 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c103
*+ bl_0_103 br_0_103 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c103
*+ bl_0_103 br_0_103 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c103
*+ bl_0_103 br_0_103 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c103
*+ bl_0_103 br_0_103 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c103
*+ bl_0_103 br_0_103 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c103
*+ bl_0_103 br_0_103 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c103
*+ bl_0_103 br_0_103 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c103
*+ bl_0_103 br_0_103 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c103
*+ bl_0_103 br_0_103 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c103
*+ bl_0_103 br_0_103 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c103
*+ bl_0_103 br_0_103 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c103
*+ bl_0_103 br_0_103 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c103
*+ bl_0_103 br_0_103 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c103
*+ bl_0_103 br_0_103 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c103
*+ bl_0_103 br_0_103 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c103
*+ bl_0_103 br_0_103 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c103
*+ bl_0_103 br_0_103 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c103
*+ bl_0_103 br_0_103 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c103
*+ bl_0_103 br_0_103 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c103
*+ bl_0_103 br_0_103 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c103
*+ bl_0_103 br_0_103 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c103
+ bl_0_103 br_0_103 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c104
+ bl_0_104 br_0_104 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c104
*+ bl_0_104 br_0_104 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c104
*+ bl_0_104 br_0_104 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c104
*+ bl_0_104 br_0_104 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c104
*+ bl_0_104 br_0_104 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c104
*+ bl_0_104 br_0_104 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c104
*+ bl_0_104 br_0_104 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c104
*+ bl_0_104 br_0_104 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c104
*+ bl_0_104 br_0_104 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c104
*+ bl_0_104 br_0_104 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c104
*+ bl_0_104 br_0_104 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c104
*+ bl_0_104 br_0_104 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c104
*+ bl_0_104 br_0_104 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c104
*+ bl_0_104 br_0_104 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c104
*+ bl_0_104 br_0_104 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c104
*+ bl_0_104 br_0_104 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c104
*+ bl_0_104 br_0_104 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c104
*+ bl_0_104 br_0_104 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c104
*+ bl_0_104 br_0_104 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c104
*+ bl_0_104 br_0_104 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c104
*+ bl_0_104 br_0_104 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c104
*+ bl_0_104 br_0_104 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c104
*+ bl_0_104 br_0_104 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c104
*+ bl_0_104 br_0_104 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c104
*+ bl_0_104 br_0_104 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c104
*+ bl_0_104 br_0_104 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c104
*+ bl_0_104 br_0_104 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c104
*+ bl_0_104 br_0_104 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c104
*+ bl_0_104 br_0_104 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c104
*+ bl_0_104 br_0_104 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c104
*+ bl_0_104 br_0_104 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c104
*+ bl_0_104 br_0_104 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c104
*+ bl_0_104 br_0_104 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c104
*+ bl_0_104 br_0_104 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c104
*+ bl_0_104 br_0_104 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c104
*+ bl_0_104 br_0_104 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c104
*+ bl_0_104 br_0_104 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c104
*+ bl_0_104 br_0_104 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c104
*+ bl_0_104 br_0_104 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c104
*+ bl_0_104 br_0_104 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c104
*+ bl_0_104 br_0_104 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c104
*+ bl_0_104 br_0_104 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c104
*+ bl_0_104 br_0_104 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c104
*+ bl_0_104 br_0_104 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c104
*+ bl_0_104 br_0_104 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c104
*+ bl_0_104 br_0_104 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c104
*+ bl_0_104 br_0_104 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c104
*+ bl_0_104 br_0_104 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c104
*+ bl_0_104 br_0_104 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c104
*+ bl_0_104 br_0_104 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c104
*+ bl_0_104 br_0_104 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c104
*+ bl_0_104 br_0_104 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c104
*+ bl_0_104 br_0_104 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c104
*+ bl_0_104 br_0_104 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c104
*+ bl_0_104 br_0_104 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c104
*+ bl_0_104 br_0_104 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c104
*+ bl_0_104 br_0_104 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c104
*+ bl_0_104 br_0_104 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c104
*+ bl_0_104 br_0_104 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c104
*+ bl_0_104 br_0_104 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c104
*+ bl_0_104 br_0_104 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c104
*+ bl_0_104 br_0_104 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c104
*+ bl_0_104 br_0_104 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c104
*+ bl_0_104 br_0_104 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c104
*+ bl_0_104 br_0_104 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c104
*+ bl_0_104 br_0_104 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c104
*+ bl_0_104 br_0_104 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c104
*+ bl_0_104 br_0_104 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c104
*+ bl_0_104 br_0_104 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c104
*+ bl_0_104 br_0_104 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c104
*+ bl_0_104 br_0_104 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c104
*+ bl_0_104 br_0_104 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c104
*+ bl_0_104 br_0_104 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c104
*+ bl_0_104 br_0_104 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c104
*+ bl_0_104 br_0_104 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c104
*+ bl_0_104 br_0_104 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c104
*+ bl_0_104 br_0_104 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c104
*+ bl_0_104 br_0_104 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c104
*+ bl_0_104 br_0_104 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c104
*+ bl_0_104 br_0_104 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c104
*+ bl_0_104 br_0_104 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c104
*+ bl_0_104 br_0_104 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c104
*+ bl_0_104 br_0_104 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c104
*+ bl_0_104 br_0_104 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c104
*+ bl_0_104 br_0_104 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c104
*+ bl_0_104 br_0_104 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c104
*+ bl_0_104 br_0_104 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c104
*+ bl_0_104 br_0_104 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c104
*+ bl_0_104 br_0_104 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c104
*+ bl_0_104 br_0_104 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c104
*+ bl_0_104 br_0_104 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c104
*+ bl_0_104 br_0_104 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c104
*+ bl_0_104 br_0_104 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c104
*+ bl_0_104 br_0_104 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c104
*+ bl_0_104 br_0_104 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c104
*+ bl_0_104 br_0_104 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c104
*+ bl_0_104 br_0_104 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c104
*+ bl_0_104 br_0_104 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c104
*+ bl_0_104 br_0_104 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c104
*+ bl_0_104 br_0_104 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c104
*+ bl_0_104 br_0_104 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c104
*+ bl_0_104 br_0_104 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c104
*+ bl_0_104 br_0_104 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c104
*+ bl_0_104 br_0_104 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c104
*+ bl_0_104 br_0_104 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c104
*+ bl_0_104 br_0_104 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c104
*+ bl_0_104 br_0_104 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c104
*+ bl_0_104 br_0_104 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c104
*+ bl_0_104 br_0_104 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c104
*+ bl_0_104 br_0_104 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c104
*+ bl_0_104 br_0_104 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c104
*+ bl_0_104 br_0_104 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c104
*+ bl_0_104 br_0_104 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c104
*+ bl_0_104 br_0_104 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c104
*+ bl_0_104 br_0_104 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c104
*+ bl_0_104 br_0_104 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c104
*+ bl_0_104 br_0_104 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c104
*+ bl_0_104 br_0_104 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c104
*+ bl_0_104 br_0_104 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c104
*+ bl_0_104 br_0_104 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c104
*+ bl_0_104 br_0_104 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c104
*+ bl_0_104 br_0_104 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c104
*+ bl_0_104 br_0_104 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c104
*+ bl_0_104 br_0_104 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c104
*+ bl_0_104 br_0_104 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c104
*+ bl_0_104 br_0_104 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c104
*+ bl_0_104 br_0_104 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c104
+ bl_0_104 br_0_104 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c105
+ bl_0_105 br_0_105 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c105
*+ bl_0_105 br_0_105 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c105
*+ bl_0_105 br_0_105 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c105
*+ bl_0_105 br_0_105 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c105
*+ bl_0_105 br_0_105 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c105
*+ bl_0_105 br_0_105 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c105
*+ bl_0_105 br_0_105 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c105
*+ bl_0_105 br_0_105 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c105
*+ bl_0_105 br_0_105 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c105
*+ bl_0_105 br_0_105 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c105
*+ bl_0_105 br_0_105 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c105
*+ bl_0_105 br_0_105 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c105
*+ bl_0_105 br_0_105 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c105
*+ bl_0_105 br_0_105 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c105
*+ bl_0_105 br_0_105 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c105
*+ bl_0_105 br_0_105 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c105
*+ bl_0_105 br_0_105 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c105
*+ bl_0_105 br_0_105 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c105
*+ bl_0_105 br_0_105 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c105
*+ bl_0_105 br_0_105 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c105
*+ bl_0_105 br_0_105 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c105
*+ bl_0_105 br_0_105 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c105
*+ bl_0_105 br_0_105 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c105
*+ bl_0_105 br_0_105 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c105
*+ bl_0_105 br_0_105 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c105
*+ bl_0_105 br_0_105 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c105
*+ bl_0_105 br_0_105 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c105
*+ bl_0_105 br_0_105 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c105
*+ bl_0_105 br_0_105 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c105
*+ bl_0_105 br_0_105 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c105
*+ bl_0_105 br_0_105 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c105
*+ bl_0_105 br_0_105 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c105
*+ bl_0_105 br_0_105 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c105
*+ bl_0_105 br_0_105 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c105
*+ bl_0_105 br_0_105 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c105
*+ bl_0_105 br_0_105 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c105
*+ bl_0_105 br_0_105 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c105
*+ bl_0_105 br_0_105 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c105
*+ bl_0_105 br_0_105 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c105
*+ bl_0_105 br_0_105 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c105
*+ bl_0_105 br_0_105 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c105
*+ bl_0_105 br_0_105 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c105
*+ bl_0_105 br_0_105 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c105
*+ bl_0_105 br_0_105 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c105
*+ bl_0_105 br_0_105 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c105
*+ bl_0_105 br_0_105 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c105
*+ bl_0_105 br_0_105 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c105
*+ bl_0_105 br_0_105 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c105
*+ bl_0_105 br_0_105 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c105
*+ bl_0_105 br_0_105 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c105
*+ bl_0_105 br_0_105 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c105
*+ bl_0_105 br_0_105 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c105
*+ bl_0_105 br_0_105 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c105
*+ bl_0_105 br_0_105 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c105
*+ bl_0_105 br_0_105 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c105
*+ bl_0_105 br_0_105 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c105
*+ bl_0_105 br_0_105 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c105
*+ bl_0_105 br_0_105 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c105
*+ bl_0_105 br_0_105 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c105
*+ bl_0_105 br_0_105 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c105
*+ bl_0_105 br_0_105 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c105
*+ bl_0_105 br_0_105 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c105
*+ bl_0_105 br_0_105 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c105
*+ bl_0_105 br_0_105 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c105
*+ bl_0_105 br_0_105 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c105
*+ bl_0_105 br_0_105 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c105
*+ bl_0_105 br_0_105 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c105
*+ bl_0_105 br_0_105 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c105
*+ bl_0_105 br_0_105 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c105
*+ bl_0_105 br_0_105 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c105
*+ bl_0_105 br_0_105 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c105
*+ bl_0_105 br_0_105 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c105
*+ bl_0_105 br_0_105 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c105
*+ bl_0_105 br_0_105 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c105
*+ bl_0_105 br_0_105 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c105
*+ bl_0_105 br_0_105 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c105
*+ bl_0_105 br_0_105 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c105
*+ bl_0_105 br_0_105 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c105
*+ bl_0_105 br_0_105 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c105
*+ bl_0_105 br_0_105 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c105
*+ bl_0_105 br_0_105 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c105
*+ bl_0_105 br_0_105 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c105
*+ bl_0_105 br_0_105 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c105
*+ bl_0_105 br_0_105 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c105
*+ bl_0_105 br_0_105 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c105
*+ bl_0_105 br_0_105 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c105
*+ bl_0_105 br_0_105 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c105
*+ bl_0_105 br_0_105 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c105
*+ bl_0_105 br_0_105 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c105
*+ bl_0_105 br_0_105 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c105
*+ bl_0_105 br_0_105 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c105
*+ bl_0_105 br_0_105 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c105
*+ bl_0_105 br_0_105 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c105
*+ bl_0_105 br_0_105 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c105
*+ bl_0_105 br_0_105 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c105
*+ bl_0_105 br_0_105 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c105
*+ bl_0_105 br_0_105 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c105
*+ bl_0_105 br_0_105 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c105
*+ bl_0_105 br_0_105 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c105
*+ bl_0_105 br_0_105 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c105
*+ bl_0_105 br_0_105 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c105
*+ bl_0_105 br_0_105 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c105
*+ bl_0_105 br_0_105 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c105
*+ bl_0_105 br_0_105 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c105
*+ bl_0_105 br_0_105 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c105
*+ bl_0_105 br_0_105 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c105
*+ bl_0_105 br_0_105 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c105
*+ bl_0_105 br_0_105 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c105
*+ bl_0_105 br_0_105 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c105
*+ bl_0_105 br_0_105 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c105
*+ bl_0_105 br_0_105 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c105
*+ bl_0_105 br_0_105 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c105
*+ bl_0_105 br_0_105 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c105
*+ bl_0_105 br_0_105 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c105
*+ bl_0_105 br_0_105 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c105
*+ bl_0_105 br_0_105 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c105
*+ bl_0_105 br_0_105 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c105
*+ bl_0_105 br_0_105 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c105
*+ bl_0_105 br_0_105 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c105
*+ bl_0_105 br_0_105 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c105
*+ bl_0_105 br_0_105 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c105
*+ bl_0_105 br_0_105 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c105
*+ bl_0_105 br_0_105 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c105
*+ bl_0_105 br_0_105 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c105
*+ bl_0_105 br_0_105 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c105
*+ bl_0_105 br_0_105 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c105
*+ bl_0_105 br_0_105 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c105
+ bl_0_105 br_0_105 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c106
+ bl_0_106 br_0_106 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c106
*+ bl_0_106 br_0_106 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c106
*+ bl_0_106 br_0_106 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c106
*+ bl_0_106 br_0_106 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c106
*+ bl_0_106 br_0_106 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c106
*+ bl_0_106 br_0_106 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c106
*+ bl_0_106 br_0_106 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c106
*+ bl_0_106 br_0_106 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c106
*+ bl_0_106 br_0_106 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c106
*+ bl_0_106 br_0_106 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c106
*+ bl_0_106 br_0_106 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c106
*+ bl_0_106 br_0_106 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c106
*+ bl_0_106 br_0_106 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c106
*+ bl_0_106 br_0_106 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c106
*+ bl_0_106 br_0_106 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c106
*+ bl_0_106 br_0_106 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c106
*+ bl_0_106 br_0_106 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c106
*+ bl_0_106 br_0_106 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c106
*+ bl_0_106 br_0_106 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c106
*+ bl_0_106 br_0_106 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c106
*+ bl_0_106 br_0_106 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c106
*+ bl_0_106 br_0_106 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c106
*+ bl_0_106 br_0_106 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c106
*+ bl_0_106 br_0_106 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c106
*+ bl_0_106 br_0_106 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c106
*+ bl_0_106 br_0_106 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c106
*+ bl_0_106 br_0_106 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c106
*+ bl_0_106 br_0_106 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c106
*+ bl_0_106 br_0_106 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c106
*+ bl_0_106 br_0_106 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c106
*+ bl_0_106 br_0_106 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c106
*+ bl_0_106 br_0_106 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c106
*+ bl_0_106 br_0_106 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c106
*+ bl_0_106 br_0_106 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c106
*+ bl_0_106 br_0_106 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c106
*+ bl_0_106 br_0_106 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c106
*+ bl_0_106 br_0_106 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c106
*+ bl_0_106 br_0_106 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c106
*+ bl_0_106 br_0_106 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c106
*+ bl_0_106 br_0_106 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c106
*+ bl_0_106 br_0_106 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c106
*+ bl_0_106 br_0_106 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c106
*+ bl_0_106 br_0_106 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c106
*+ bl_0_106 br_0_106 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c106
*+ bl_0_106 br_0_106 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c106
*+ bl_0_106 br_0_106 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c106
*+ bl_0_106 br_0_106 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c106
*+ bl_0_106 br_0_106 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c106
*+ bl_0_106 br_0_106 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c106
*+ bl_0_106 br_0_106 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c106
*+ bl_0_106 br_0_106 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c106
*+ bl_0_106 br_0_106 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c106
*+ bl_0_106 br_0_106 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c106
*+ bl_0_106 br_0_106 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c106
*+ bl_0_106 br_0_106 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c106
*+ bl_0_106 br_0_106 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c106
*+ bl_0_106 br_0_106 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c106
*+ bl_0_106 br_0_106 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c106
*+ bl_0_106 br_0_106 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c106
*+ bl_0_106 br_0_106 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c106
*+ bl_0_106 br_0_106 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c106
*+ bl_0_106 br_0_106 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c106
*+ bl_0_106 br_0_106 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c106
*+ bl_0_106 br_0_106 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c106
*+ bl_0_106 br_0_106 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c106
*+ bl_0_106 br_0_106 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c106
*+ bl_0_106 br_0_106 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c106
*+ bl_0_106 br_0_106 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c106
*+ bl_0_106 br_0_106 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c106
*+ bl_0_106 br_0_106 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c106
*+ bl_0_106 br_0_106 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c106
*+ bl_0_106 br_0_106 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c106
*+ bl_0_106 br_0_106 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c106
*+ bl_0_106 br_0_106 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c106
*+ bl_0_106 br_0_106 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c106
*+ bl_0_106 br_0_106 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c106
*+ bl_0_106 br_0_106 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c106
*+ bl_0_106 br_0_106 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c106
*+ bl_0_106 br_0_106 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c106
*+ bl_0_106 br_0_106 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c106
*+ bl_0_106 br_0_106 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c106
*+ bl_0_106 br_0_106 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c106
*+ bl_0_106 br_0_106 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c106
*+ bl_0_106 br_0_106 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c106
*+ bl_0_106 br_0_106 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c106
*+ bl_0_106 br_0_106 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c106
*+ bl_0_106 br_0_106 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c106
*+ bl_0_106 br_0_106 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c106
*+ bl_0_106 br_0_106 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c106
*+ bl_0_106 br_0_106 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c106
*+ bl_0_106 br_0_106 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c106
*+ bl_0_106 br_0_106 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c106
*+ bl_0_106 br_0_106 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c106
*+ bl_0_106 br_0_106 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c106
*+ bl_0_106 br_0_106 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c106
*+ bl_0_106 br_0_106 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c106
*+ bl_0_106 br_0_106 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c106
*+ bl_0_106 br_0_106 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c106
*+ bl_0_106 br_0_106 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c106
*+ bl_0_106 br_0_106 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c106
*+ bl_0_106 br_0_106 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c106
*+ bl_0_106 br_0_106 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c106
*+ bl_0_106 br_0_106 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c106
*+ bl_0_106 br_0_106 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c106
*+ bl_0_106 br_0_106 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c106
*+ bl_0_106 br_0_106 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c106
*+ bl_0_106 br_0_106 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c106
*+ bl_0_106 br_0_106 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c106
*+ bl_0_106 br_0_106 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c106
*+ bl_0_106 br_0_106 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c106
*+ bl_0_106 br_0_106 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c106
*+ bl_0_106 br_0_106 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c106
*+ bl_0_106 br_0_106 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c106
*+ bl_0_106 br_0_106 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c106
*+ bl_0_106 br_0_106 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c106
*+ bl_0_106 br_0_106 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c106
*+ bl_0_106 br_0_106 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c106
*+ bl_0_106 br_0_106 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c106
*+ bl_0_106 br_0_106 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c106
*+ bl_0_106 br_0_106 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c106
*+ bl_0_106 br_0_106 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c106
*+ bl_0_106 br_0_106 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c106
*+ bl_0_106 br_0_106 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c106
*+ bl_0_106 br_0_106 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c106
*+ bl_0_106 br_0_106 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c106
*+ bl_0_106 br_0_106 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c106
*+ bl_0_106 br_0_106 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c106
+ bl_0_106 br_0_106 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c107
+ bl_0_107 br_0_107 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c107
*+ bl_0_107 br_0_107 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c107
*+ bl_0_107 br_0_107 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c107
*+ bl_0_107 br_0_107 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c107
*+ bl_0_107 br_0_107 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c107
*+ bl_0_107 br_0_107 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c107
*+ bl_0_107 br_0_107 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c107
*+ bl_0_107 br_0_107 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c107
*+ bl_0_107 br_0_107 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c107
*+ bl_0_107 br_0_107 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c107
*+ bl_0_107 br_0_107 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c107
*+ bl_0_107 br_0_107 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c107
*+ bl_0_107 br_0_107 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c107
*+ bl_0_107 br_0_107 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c107
*+ bl_0_107 br_0_107 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c107
*+ bl_0_107 br_0_107 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c107
*+ bl_0_107 br_0_107 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c107
*+ bl_0_107 br_0_107 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c107
*+ bl_0_107 br_0_107 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c107
*+ bl_0_107 br_0_107 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c107
*+ bl_0_107 br_0_107 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c107
*+ bl_0_107 br_0_107 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c107
*+ bl_0_107 br_0_107 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c107
*+ bl_0_107 br_0_107 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c107
*+ bl_0_107 br_0_107 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c107
*+ bl_0_107 br_0_107 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c107
*+ bl_0_107 br_0_107 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c107
*+ bl_0_107 br_0_107 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c107
*+ bl_0_107 br_0_107 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c107
*+ bl_0_107 br_0_107 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c107
*+ bl_0_107 br_0_107 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c107
*+ bl_0_107 br_0_107 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c107
*+ bl_0_107 br_0_107 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c107
*+ bl_0_107 br_0_107 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c107
*+ bl_0_107 br_0_107 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c107
*+ bl_0_107 br_0_107 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c107
*+ bl_0_107 br_0_107 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c107
*+ bl_0_107 br_0_107 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c107
*+ bl_0_107 br_0_107 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c107
*+ bl_0_107 br_0_107 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c107
*+ bl_0_107 br_0_107 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c107
*+ bl_0_107 br_0_107 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c107
*+ bl_0_107 br_0_107 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c107
*+ bl_0_107 br_0_107 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c107
*+ bl_0_107 br_0_107 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c107
*+ bl_0_107 br_0_107 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c107
*+ bl_0_107 br_0_107 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c107
*+ bl_0_107 br_0_107 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c107
*+ bl_0_107 br_0_107 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c107
*+ bl_0_107 br_0_107 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c107
*+ bl_0_107 br_0_107 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c107
*+ bl_0_107 br_0_107 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c107
*+ bl_0_107 br_0_107 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c107
*+ bl_0_107 br_0_107 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c107
*+ bl_0_107 br_0_107 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c107
*+ bl_0_107 br_0_107 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c107
*+ bl_0_107 br_0_107 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c107
*+ bl_0_107 br_0_107 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c107
*+ bl_0_107 br_0_107 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c107
*+ bl_0_107 br_0_107 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c107
*+ bl_0_107 br_0_107 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c107
*+ bl_0_107 br_0_107 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c107
*+ bl_0_107 br_0_107 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c107
*+ bl_0_107 br_0_107 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c107
*+ bl_0_107 br_0_107 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c107
*+ bl_0_107 br_0_107 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c107
*+ bl_0_107 br_0_107 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c107
*+ bl_0_107 br_0_107 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c107
*+ bl_0_107 br_0_107 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c107
*+ bl_0_107 br_0_107 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c107
*+ bl_0_107 br_0_107 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c107
*+ bl_0_107 br_0_107 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c107
*+ bl_0_107 br_0_107 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c107
*+ bl_0_107 br_0_107 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c107
*+ bl_0_107 br_0_107 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c107
*+ bl_0_107 br_0_107 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c107
*+ bl_0_107 br_0_107 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c107
*+ bl_0_107 br_0_107 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c107
*+ bl_0_107 br_0_107 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c107
*+ bl_0_107 br_0_107 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c107
*+ bl_0_107 br_0_107 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c107
*+ bl_0_107 br_0_107 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c107
*+ bl_0_107 br_0_107 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c107
*+ bl_0_107 br_0_107 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c107
*+ bl_0_107 br_0_107 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c107
*+ bl_0_107 br_0_107 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c107
*+ bl_0_107 br_0_107 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c107
*+ bl_0_107 br_0_107 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c107
*+ bl_0_107 br_0_107 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c107
*+ bl_0_107 br_0_107 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c107
*+ bl_0_107 br_0_107 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c107
*+ bl_0_107 br_0_107 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c107
*+ bl_0_107 br_0_107 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c107
*+ bl_0_107 br_0_107 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c107
*+ bl_0_107 br_0_107 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c107
*+ bl_0_107 br_0_107 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c107
*+ bl_0_107 br_0_107 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c107
*+ bl_0_107 br_0_107 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c107
*+ bl_0_107 br_0_107 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c107
*+ bl_0_107 br_0_107 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c107
*+ bl_0_107 br_0_107 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c107
*+ bl_0_107 br_0_107 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c107
*+ bl_0_107 br_0_107 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c107
*+ bl_0_107 br_0_107 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c107
*+ bl_0_107 br_0_107 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c107
*+ bl_0_107 br_0_107 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c107
*+ bl_0_107 br_0_107 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c107
*+ bl_0_107 br_0_107 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c107
*+ bl_0_107 br_0_107 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c107
*+ bl_0_107 br_0_107 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c107
*+ bl_0_107 br_0_107 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c107
*+ bl_0_107 br_0_107 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c107
*+ bl_0_107 br_0_107 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c107
*+ bl_0_107 br_0_107 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c107
*+ bl_0_107 br_0_107 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c107
*+ bl_0_107 br_0_107 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c107
*+ bl_0_107 br_0_107 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c107
*+ bl_0_107 br_0_107 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c107
*+ bl_0_107 br_0_107 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c107
*+ bl_0_107 br_0_107 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c107
*+ bl_0_107 br_0_107 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c107
*+ bl_0_107 br_0_107 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c107
*+ bl_0_107 br_0_107 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c107
*+ bl_0_107 br_0_107 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c107
*+ bl_0_107 br_0_107 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c107
*+ bl_0_107 br_0_107 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c107
*+ bl_0_107 br_0_107 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c107
+ bl_0_107 br_0_107 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c108
+ bl_0_108 br_0_108 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c108
*+ bl_0_108 br_0_108 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c108
*+ bl_0_108 br_0_108 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c108
*+ bl_0_108 br_0_108 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c108
*+ bl_0_108 br_0_108 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c108
*+ bl_0_108 br_0_108 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c108
*+ bl_0_108 br_0_108 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c108
*+ bl_0_108 br_0_108 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c108
*+ bl_0_108 br_0_108 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c108
*+ bl_0_108 br_0_108 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c108
*+ bl_0_108 br_0_108 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c108
*+ bl_0_108 br_0_108 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c108
*+ bl_0_108 br_0_108 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c108
*+ bl_0_108 br_0_108 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c108
*+ bl_0_108 br_0_108 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c108
*+ bl_0_108 br_0_108 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c108
*+ bl_0_108 br_0_108 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c108
*+ bl_0_108 br_0_108 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c108
*+ bl_0_108 br_0_108 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c108
*+ bl_0_108 br_0_108 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c108
*+ bl_0_108 br_0_108 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c108
*+ bl_0_108 br_0_108 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c108
*+ bl_0_108 br_0_108 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c108
*+ bl_0_108 br_0_108 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c108
*+ bl_0_108 br_0_108 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c108
*+ bl_0_108 br_0_108 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c108
*+ bl_0_108 br_0_108 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c108
*+ bl_0_108 br_0_108 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c108
*+ bl_0_108 br_0_108 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c108
*+ bl_0_108 br_0_108 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c108
*+ bl_0_108 br_0_108 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c108
*+ bl_0_108 br_0_108 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c108
*+ bl_0_108 br_0_108 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c108
*+ bl_0_108 br_0_108 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c108
*+ bl_0_108 br_0_108 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c108
*+ bl_0_108 br_0_108 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c108
*+ bl_0_108 br_0_108 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c108
*+ bl_0_108 br_0_108 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c108
*+ bl_0_108 br_0_108 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c108
*+ bl_0_108 br_0_108 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c108
*+ bl_0_108 br_0_108 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c108
*+ bl_0_108 br_0_108 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c108
*+ bl_0_108 br_0_108 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c108
*+ bl_0_108 br_0_108 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c108
*+ bl_0_108 br_0_108 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c108
*+ bl_0_108 br_0_108 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c108
*+ bl_0_108 br_0_108 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c108
*+ bl_0_108 br_0_108 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c108
*+ bl_0_108 br_0_108 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c108
*+ bl_0_108 br_0_108 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c108
*+ bl_0_108 br_0_108 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c108
*+ bl_0_108 br_0_108 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c108
*+ bl_0_108 br_0_108 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c108
*+ bl_0_108 br_0_108 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c108
*+ bl_0_108 br_0_108 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c108
*+ bl_0_108 br_0_108 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c108
*+ bl_0_108 br_0_108 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c108
*+ bl_0_108 br_0_108 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c108
*+ bl_0_108 br_0_108 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c108
*+ bl_0_108 br_0_108 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c108
*+ bl_0_108 br_0_108 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c108
*+ bl_0_108 br_0_108 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c108
*+ bl_0_108 br_0_108 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c108
*+ bl_0_108 br_0_108 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c108
*+ bl_0_108 br_0_108 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c108
*+ bl_0_108 br_0_108 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c108
*+ bl_0_108 br_0_108 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c108
*+ bl_0_108 br_0_108 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c108
*+ bl_0_108 br_0_108 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c108
*+ bl_0_108 br_0_108 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c108
*+ bl_0_108 br_0_108 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c108
*+ bl_0_108 br_0_108 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c108
*+ bl_0_108 br_0_108 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c108
*+ bl_0_108 br_0_108 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c108
*+ bl_0_108 br_0_108 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c108
*+ bl_0_108 br_0_108 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c108
*+ bl_0_108 br_0_108 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c108
*+ bl_0_108 br_0_108 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c108
*+ bl_0_108 br_0_108 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c108
*+ bl_0_108 br_0_108 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c108
*+ bl_0_108 br_0_108 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c108
*+ bl_0_108 br_0_108 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c108
*+ bl_0_108 br_0_108 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c108
*+ bl_0_108 br_0_108 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c108
*+ bl_0_108 br_0_108 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c108
*+ bl_0_108 br_0_108 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c108
*+ bl_0_108 br_0_108 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c108
*+ bl_0_108 br_0_108 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c108
*+ bl_0_108 br_0_108 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c108
*+ bl_0_108 br_0_108 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c108
*+ bl_0_108 br_0_108 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c108
*+ bl_0_108 br_0_108 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c108
*+ bl_0_108 br_0_108 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c108
*+ bl_0_108 br_0_108 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c108
*+ bl_0_108 br_0_108 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c108
*+ bl_0_108 br_0_108 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c108
*+ bl_0_108 br_0_108 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c108
*+ bl_0_108 br_0_108 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c108
*+ bl_0_108 br_0_108 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c108
*+ bl_0_108 br_0_108 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c108
*+ bl_0_108 br_0_108 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c108
*+ bl_0_108 br_0_108 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c108
*+ bl_0_108 br_0_108 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c108
*+ bl_0_108 br_0_108 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c108
*+ bl_0_108 br_0_108 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c108
*+ bl_0_108 br_0_108 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c108
*+ bl_0_108 br_0_108 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c108
*+ bl_0_108 br_0_108 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c108
*+ bl_0_108 br_0_108 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c108
*+ bl_0_108 br_0_108 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c108
*+ bl_0_108 br_0_108 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c108
*+ bl_0_108 br_0_108 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c108
*+ bl_0_108 br_0_108 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c108
*+ bl_0_108 br_0_108 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c108
*+ bl_0_108 br_0_108 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c108
*+ bl_0_108 br_0_108 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c108
*+ bl_0_108 br_0_108 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c108
*+ bl_0_108 br_0_108 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c108
*+ bl_0_108 br_0_108 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c108
*+ bl_0_108 br_0_108 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c108
*+ bl_0_108 br_0_108 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c108
*+ bl_0_108 br_0_108 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c108
*+ bl_0_108 br_0_108 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c108
*+ bl_0_108 br_0_108 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c108
*+ bl_0_108 br_0_108 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c108
*+ bl_0_108 br_0_108 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c108
*+ bl_0_108 br_0_108 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c108
+ bl_0_108 br_0_108 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c109
+ bl_0_109 br_0_109 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c109
*+ bl_0_109 br_0_109 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c109
*+ bl_0_109 br_0_109 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c109
*+ bl_0_109 br_0_109 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c109
*+ bl_0_109 br_0_109 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c109
*+ bl_0_109 br_0_109 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c109
*+ bl_0_109 br_0_109 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c109
*+ bl_0_109 br_0_109 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c109
*+ bl_0_109 br_0_109 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c109
*+ bl_0_109 br_0_109 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c109
*+ bl_0_109 br_0_109 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c109
*+ bl_0_109 br_0_109 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c109
*+ bl_0_109 br_0_109 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c109
*+ bl_0_109 br_0_109 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c109
*+ bl_0_109 br_0_109 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c109
*+ bl_0_109 br_0_109 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c109
*+ bl_0_109 br_0_109 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c109
*+ bl_0_109 br_0_109 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c109
*+ bl_0_109 br_0_109 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c109
*+ bl_0_109 br_0_109 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c109
*+ bl_0_109 br_0_109 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c109
*+ bl_0_109 br_0_109 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c109
*+ bl_0_109 br_0_109 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c109
*+ bl_0_109 br_0_109 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c109
*+ bl_0_109 br_0_109 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c109
*+ bl_0_109 br_0_109 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c109
*+ bl_0_109 br_0_109 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c109
*+ bl_0_109 br_0_109 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c109
*+ bl_0_109 br_0_109 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c109
*+ bl_0_109 br_0_109 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c109
*+ bl_0_109 br_0_109 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c109
*+ bl_0_109 br_0_109 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c109
*+ bl_0_109 br_0_109 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c109
*+ bl_0_109 br_0_109 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c109
*+ bl_0_109 br_0_109 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c109
*+ bl_0_109 br_0_109 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c109
*+ bl_0_109 br_0_109 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c109
*+ bl_0_109 br_0_109 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c109
*+ bl_0_109 br_0_109 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c109
*+ bl_0_109 br_0_109 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c109
*+ bl_0_109 br_0_109 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c109
*+ bl_0_109 br_0_109 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c109
*+ bl_0_109 br_0_109 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c109
*+ bl_0_109 br_0_109 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c109
*+ bl_0_109 br_0_109 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c109
*+ bl_0_109 br_0_109 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c109
*+ bl_0_109 br_0_109 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c109
*+ bl_0_109 br_0_109 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c109
*+ bl_0_109 br_0_109 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c109
*+ bl_0_109 br_0_109 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c109
*+ bl_0_109 br_0_109 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c109
*+ bl_0_109 br_0_109 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c109
*+ bl_0_109 br_0_109 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c109
*+ bl_0_109 br_0_109 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c109
*+ bl_0_109 br_0_109 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c109
*+ bl_0_109 br_0_109 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c109
*+ bl_0_109 br_0_109 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c109
*+ bl_0_109 br_0_109 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c109
*+ bl_0_109 br_0_109 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c109
*+ bl_0_109 br_0_109 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c109
*+ bl_0_109 br_0_109 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c109
*+ bl_0_109 br_0_109 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c109
*+ bl_0_109 br_0_109 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c109
*+ bl_0_109 br_0_109 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c109
*+ bl_0_109 br_0_109 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c109
*+ bl_0_109 br_0_109 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c109
*+ bl_0_109 br_0_109 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c109
*+ bl_0_109 br_0_109 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c109
*+ bl_0_109 br_0_109 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c109
*+ bl_0_109 br_0_109 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c109
*+ bl_0_109 br_0_109 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c109
*+ bl_0_109 br_0_109 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c109
*+ bl_0_109 br_0_109 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c109
*+ bl_0_109 br_0_109 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c109
*+ bl_0_109 br_0_109 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c109
*+ bl_0_109 br_0_109 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c109
*+ bl_0_109 br_0_109 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c109
*+ bl_0_109 br_0_109 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c109
*+ bl_0_109 br_0_109 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c109
*+ bl_0_109 br_0_109 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c109
*+ bl_0_109 br_0_109 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c109
*+ bl_0_109 br_0_109 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c109
*+ bl_0_109 br_0_109 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c109
*+ bl_0_109 br_0_109 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c109
*+ bl_0_109 br_0_109 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c109
*+ bl_0_109 br_0_109 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c109
*+ bl_0_109 br_0_109 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c109
*+ bl_0_109 br_0_109 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c109
*+ bl_0_109 br_0_109 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c109
*+ bl_0_109 br_0_109 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c109
*+ bl_0_109 br_0_109 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c109
*+ bl_0_109 br_0_109 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c109
*+ bl_0_109 br_0_109 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c109
*+ bl_0_109 br_0_109 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c109
*+ bl_0_109 br_0_109 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c109
*+ bl_0_109 br_0_109 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c109
*+ bl_0_109 br_0_109 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c109
*+ bl_0_109 br_0_109 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c109
*+ bl_0_109 br_0_109 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c109
*+ bl_0_109 br_0_109 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c109
*+ bl_0_109 br_0_109 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c109
*+ bl_0_109 br_0_109 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c109
*+ bl_0_109 br_0_109 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c109
*+ bl_0_109 br_0_109 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c109
*+ bl_0_109 br_0_109 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c109
*+ bl_0_109 br_0_109 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c109
*+ bl_0_109 br_0_109 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c109
*+ bl_0_109 br_0_109 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c109
*+ bl_0_109 br_0_109 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c109
*+ bl_0_109 br_0_109 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c109
*+ bl_0_109 br_0_109 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c109
*+ bl_0_109 br_0_109 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c109
*+ bl_0_109 br_0_109 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c109
*+ bl_0_109 br_0_109 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c109
*+ bl_0_109 br_0_109 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c109
*+ bl_0_109 br_0_109 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c109
*+ bl_0_109 br_0_109 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c109
*+ bl_0_109 br_0_109 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c109
*+ bl_0_109 br_0_109 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c109
*+ bl_0_109 br_0_109 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c109
*+ bl_0_109 br_0_109 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c109
*+ bl_0_109 br_0_109 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c109
*+ bl_0_109 br_0_109 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c109
*+ bl_0_109 br_0_109 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c109
*+ bl_0_109 br_0_109 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c109
*+ bl_0_109 br_0_109 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c109
*+ bl_0_109 br_0_109 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c109
+ bl_0_109 br_0_109 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c110
+ bl_0_110 br_0_110 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c110
*+ bl_0_110 br_0_110 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c110
*+ bl_0_110 br_0_110 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c110
*+ bl_0_110 br_0_110 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c110
*+ bl_0_110 br_0_110 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c110
*+ bl_0_110 br_0_110 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c110
*+ bl_0_110 br_0_110 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c110
*+ bl_0_110 br_0_110 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c110
*+ bl_0_110 br_0_110 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c110
*+ bl_0_110 br_0_110 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c110
*+ bl_0_110 br_0_110 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c110
*+ bl_0_110 br_0_110 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c110
*+ bl_0_110 br_0_110 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c110
*+ bl_0_110 br_0_110 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c110
*+ bl_0_110 br_0_110 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c110
*+ bl_0_110 br_0_110 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c110
*+ bl_0_110 br_0_110 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c110
*+ bl_0_110 br_0_110 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c110
*+ bl_0_110 br_0_110 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c110
*+ bl_0_110 br_0_110 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c110
*+ bl_0_110 br_0_110 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c110
*+ bl_0_110 br_0_110 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c110
*+ bl_0_110 br_0_110 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c110
*+ bl_0_110 br_0_110 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c110
*+ bl_0_110 br_0_110 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c110
*+ bl_0_110 br_0_110 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c110
*+ bl_0_110 br_0_110 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c110
*+ bl_0_110 br_0_110 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c110
*+ bl_0_110 br_0_110 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c110
*+ bl_0_110 br_0_110 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c110
*+ bl_0_110 br_0_110 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c110
*+ bl_0_110 br_0_110 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c110
*+ bl_0_110 br_0_110 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c110
*+ bl_0_110 br_0_110 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c110
*+ bl_0_110 br_0_110 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c110
*+ bl_0_110 br_0_110 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c110
*+ bl_0_110 br_0_110 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c110
*+ bl_0_110 br_0_110 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c110
*+ bl_0_110 br_0_110 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c110
*+ bl_0_110 br_0_110 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c110
*+ bl_0_110 br_0_110 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c110
*+ bl_0_110 br_0_110 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c110
*+ bl_0_110 br_0_110 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c110
*+ bl_0_110 br_0_110 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c110
*+ bl_0_110 br_0_110 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c110
*+ bl_0_110 br_0_110 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c110
*+ bl_0_110 br_0_110 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c110
*+ bl_0_110 br_0_110 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c110
*+ bl_0_110 br_0_110 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c110
*+ bl_0_110 br_0_110 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c110
*+ bl_0_110 br_0_110 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c110
*+ bl_0_110 br_0_110 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c110
*+ bl_0_110 br_0_110 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c110
*+ bl_0_110 br_0_110 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c110
*+ bl_0_110 br_0_110 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c110
*+ bl_0_110 br_0_110 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c110
*+ bl_0_110 br_0_110 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c110
*+ bl_0_110 br_0_110 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c110
*+ bl_0_110 br_0_110 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c110
*+ bl_0_110 br_0_110 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c110
*+ bl_0_110 br_0_110 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c110
*+ bl_0_110 br_0_110 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c110
*+ bl_0_110 br_0_110 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c110
*+ bl_0_110 br_0_110 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c110
*+ bl_0_110 br_0_110 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c110
*+ bl_0_110 br_0_110 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c110
*+ bl_0_110 br_0_110 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c110
*+ bl_0_110 br_0_110 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c110
*+ bl_0_110 br_0_110 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c110
*+ bl_0_110 br_0_110 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c110
*+ bl_0_110 br_0_110 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c110
*+ bl_0_110 br_0_110 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c110
*+ bl_0_110 br_0_110 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c110
*+ bl_0_110 br_0_110 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c110
*+ bl_0_110 br_0_110 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c110
*+ bl_0_110 br_0_110 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c110
*+ bl_0_110 br_0_110 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c110
*+ bl_0_110 br_0_110 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c110
*+ bl_0_110 br_0_110 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c110
*+ bl_0_110 br_0_110 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c110
*+ bl_0_110 br_0_110 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c110
*+ bl_0_110 br_0_110 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c110
*+ bl_0_110 br_0_110 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c110
*+ bl_0_110 br_0_110 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c110
*+ bl_0_110 br_0_110 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c110
*+ bl_0_110 br_0_110 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c110
*+ bl_0_110 br_0_110 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c110
*+ bl_0_110 br_0_110 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c110
*+ bl_0_110 br_0_110 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c110
*+ bl_0_110 br_0_110 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c110
*+ bl_0_110 br_0_110 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c110
*+ bl_0_110 br_0_110 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c110
*+ bl_0_110 br_0_110 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c110
*+ bl_0_110 br_0_110 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c110
*+ bl_0_110 br_0_110 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c110
*+ bl_0_110 br_0_110 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c110
*+ bl_0_110 br_0_110 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c110
*+ bl_0_110 br_0_110 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c110
*+ bl_0_110 br_0_110 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c110
*+ bl_0_110 br_0_110 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c110
*+ bl_0_110 br_0_110 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c110
*+ bl_0_110 br_0_110 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c110
*+ bl_0_110 br_0_110 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c110
*+ bl_0_110 br_0_110 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c110
*+ bl_0_110 br_0_110 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c110
*+ bl_0_110 br_0_110 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c110
*+ bl_0_110 br_0_110 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c110
*+ bl_0_110 br_0_110 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c110
*+ bl_0_110 br_0_110 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c110
*+ bl_0_110 br_0_110 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c110
*+ bl_0_110 br_0_110 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c110
*+ bl_0_110 br_0_110 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c110
*+ bl_0_110 br_0_110 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c110
*+ bl_0_110 br_0_110 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c110
*+ bl_0_110 br_0_110 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c110
*+ bl_0_110 br_0_110 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c110
*+ bl_0_110 br_0_110 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c110
*+ bl_0_110 br_0_110 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c110
*+ bl_0_110 br_0_110 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c110
*+ bl_0_110 br_0_110 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c110
*+ bl_0_110 br_0_110 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c110
*+ bl_0_110 br_0_110 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c110
*+ bl_0_110 br_0_110 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c110
*+ bl_0_110 br_0_110 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c110
*+ bl_0_110 br_0_110 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c110
*+ bl_0_110 br_0_110 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c110
*+ bl_0_110 br_0_110 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c110
+ bl_0_110 br_0_110 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c111
+ bl_0_111 br_0_111 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c111
*+ bl_0_111 br_0_111 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c111
*+ bl_0_111 br_0_111 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c111
*+ bl_0_111 br_0_111 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c111
*+ bl_0_111 br_0_111 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c111
*+ bl_0_111 br_0_111 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c111
*+ bl_0_111 br_0_111 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c111
*+ bl_0_111 br_0_111 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c111
*+ bl_0_111 br_0_111 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c111
*+ bl_0_111 br_0_111 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c111
*+ bl_0_111 br_0_111 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c111
*+ bl_0_111 br_0_111 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c111
*+ bl_0_111 br_0_111 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c111
*+ bl_0_111 br_0_111 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c111
*+ bl_0_111 br_0_111 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c111
*+ bl_0_111 br_0_111 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c111
*+ bl_0_111 br_0_111 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c111
*+ bl_0_111 br_0_111 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c111
*+ bl_0_111 br_0_111 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c111
*+ bl_0_111 br_0_111 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c111
*+ bl_0_111 br_0_111 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c111
*+ bl_0_111 br_0_111 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c111
*+ bl_0_111 br_0_111 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c111
*+ bl_0_111 br_0_111 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c111
*+ bl_0_111 br_0_111 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c111
*+ bl_0_111 br_0_111 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c111
*+ bl_0_111 br_0_111 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c111
*+ bl_0_111 br_0_111 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c111
*+ bl_0_111 br_0_111 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c111
*+ bl_0_111 br_0_111 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c111
*+ bl_0_111 br_0_111 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c111
*+ bl_0_111 br_0_111 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c111
*+ bl_0_111 br_0_111 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c111
*+ bl_0_111 br_0_111 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c111
*+ bl_0_111 br_0_111 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c111
*+ bl_0_111 br_0_111 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c111
*+ bl_0_111 br_0_111 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c111
*+ bl_0_111 br_0_111 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c111
*+ bl_0_111 br_0_111 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c111
*+ bl_0_111 br_0_111 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c111
*+ bl_0_111 br_0_111 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c111
*+ bl_0_111 br_0_111 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c111
*+ bl_0_111 br_0_111 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c111
*+ bl_0_111 br_0_111 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c111
*+ bl_0_111 br_0_111 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c111
*+ bl_0_111 br_0_111 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c111
*+ bl_0_111 br_0_111 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c111
*+ bl_0_111 br_0_111 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c111
*+ bl_0_111 br_0_111 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c111
*+ bl_0_111 br_0_111 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c111
*+ bl_0_111 br_0_111 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c111
*+ bl_0_111 br_0_111 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c111
*+ bl_0_111 br_0_111 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c111
*+ bl_0_111 br_0_111 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c111
*+ bl_0_111 br_0_111 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c111
*+ bl_0_111 br_0_111 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c111
*+ bl_0_111 br_0_111 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c111
*+ bl_0_111 br_0_111 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c111
*+ bl_0_111 br_0_111 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c111
*+ bl_0_111 br_0_111 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c111
*+ bl_0_111 br_0_111 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c111
*+ bl_0_111 br_0_111 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c111
*+ bl_0_111 br_0_111 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c111
*+ bl_0_111 br_0_111 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c111
*+ bl_0_111 br_0_111 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c111
*+ bl_0_111 br_0_111 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c111
*+ bl_0_111 br_0_111 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c111
*+ bl_0_111 br_0_111 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c111
*+ bl_0_111 br_0_111 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c111
*+ bl_0_111 br_0_111 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c111
*+ bl_0_111 br_0_111 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c111
*+ bl_0_111 br_0_111 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c111
*+ bl_0_111 br_0_111 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c111
*+ bl_0_111 br_0_111 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c111
*+ bl_0_111 br_0_111 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c111
*+ bl_0_111 br_0_111 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c111
*+ bl_0_111 br_0_111 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c111
*+ bl_0_111 br_0_111 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c111
*+ bl_0_111 br_0_111 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c111
*+ bl_0_111 br_0_111 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c111
*+ bl_0_111 br_0_111 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c111
*+ bl_0_111 br_0_111 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c111
*+ bl_0_111 br_0_111 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c111
*+ bl_0_111 br_0_111 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c111
*+ bl_0_111 br_0_111 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c111
*+ bl_0_111 br_0_111 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c111
*+ bl_0_111 br_0_111 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c111
*+ bl_0_111 br_0_111 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c111
*+ bl_0_111 br_0_111 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c111
*+ bl_0_111 br_0_111 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c111
*+ bl_0_111 br_0_111 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c111
*+ bl_0_111 br_0_111 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c111
*+ bl_0_111 br_0_111 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c111
*+ bl_0_111 br_0_111 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c111
*+ bl_0_111 br_0_111 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c111
*+ bl_0_111 br_0_111 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c111
*+ bl_0_111 br_0_111 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c111
*+ bl_0_111 br_0_111 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c111
*+ bl_0_111 br_0_111 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c111
*+ bl_0_111 br_0_111 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c111
*+ bl_0_111 br_0_111 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c111
*+ bl_0_111 br_0_111 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c111
*+ bl_0_111 br_0_111 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c111
*+ bl_0_111 br_0_111 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c111
*+ bl_0_111 br_0_111 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c111
*+ bl_0_111 br_0_111 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c111
*+ bl_0_111 br_0_111 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c111
*+ bl_0_111 br_0_111 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c111
*+ bl_0_111 br_0_111 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c111
*+ bl_0_111 br_0_111 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c111
*+ bl_0_111 br_0_111 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c111
*+ bl_0_111 br_0_111 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c111
*+ bl_0_111 br_0_111 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c111
*+ bl_0_111 br_0_111 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c111
*+ bl_0_111 br_0_111 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c111
*+ bl_0_111 br_0_111 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c111
*+ bl_0_111 br_0_111 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c111
*+ bl_0_111 br_0_111 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c111
*+ bl_0_111 br_0_111 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c111
*+ bl_0_111 br_0_111 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c111
*+ bl_0_111 br_0_111 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c111
*+ bl_0_111 br_0_111 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c111
*+ bl_0_111 br_0_111 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c111
*+ bl_0_111 br_0_111 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c111
*+ bl_0_111 br_0_111 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c111
*+ bl_0_111 br_0_111 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c111
*+ bl_0_111 br_0_111 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c111
+ bl_0_111 br_0_111 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c112
+ bl_0_112 br_0_112 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c112
*+ bl_0_112 br_0_112 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c112
*+ bl_0_112 br_0_112 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c112
*+ bl_0_112 br_0_112 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c112
*+ bl_0_112 br_0_112 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c112
*+ bl_0_112 br_0_112 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c112
*+ bl_0_112 br_0_112 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c112
*+ bl_0_112 br_0_112 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c112
*+ bl_0_112 br_0_112 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c112
*+ bl_0_112 br_0_112 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c112
*+ bl_0_112 br_0_112 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c112
*+ bl_0_112 br_0_112 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c112
*+ bl_0_112 br_0_112 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c112
*+ bl_0_112 br_0_112 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c112
*+ bl_0_112 br_0_112 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c112
*+ bl_0_112 br_0_112 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c112
*+ bl_0_112 br_0_112 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c112
*+ bl_0_112 br_0_112 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c112
*+ bl_0_112 br_0_112 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c112
*+ bl_0_112 br_0_112 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c112
*+ bl_0_112 br_0_112 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c112
*+ bl_0_112 br_0_112 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c112
*+ bl_0_112 br_0_112 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c112
*+ bl_0_112 br_0_112 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c112
*+ bl_0_112 br_0_112 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c112
*+ bl_0_112 br_0_112 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c112
*+ bl_0_112 br_0_112 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c112
*+ bl_0_112 br_0_112 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c112
*+ bl_0_112 br_0_112 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c112
*+ bl_0_112 br_0_112 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c112
*+ bl_0_112 br_0_112 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c112
*+ bl_0_112 br_0_112 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c112
*+ bl_0_112 br_0_112 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c112
*+ bl_0_112 br_0_112 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c112
*+ bl_0_112 br_0_112 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c112
*+ bl_0_112 br_0_112 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c112
*+ bl_0_112 br_0_112 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c112
*+ bl_0_112 br_0_112 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c112
*+ bl_0_112 br_0_112 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c112
*+ bl_0_112 br_0_112 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c112
*+ bl_0_112 br_0_112 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c112
*+ bl_0_112 br_0_112 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c112
*+ bl_0_112 br_0_112 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c112
*+ bl_0_112 br_0_112 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c112
*+ bl_0_112 br_0_112 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c112
*+ bl_0_112 br_0_112 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c112
*+ bl_0_112 br_0_112 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c112
*+ bl_0_112 br_0_112 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c112
*+ bl_0_112 br_0_112 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c112
*+ bl_0_112 br_0_112 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c112
*+ bl_0_112 br_0_112 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c112
*+ bl_0_112 br_0_112 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c112
*+ bl_0_112 br_0_112 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c112
*+ bl_0_112 br_0_112 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c112
*+ bl_0_112 br_0_112 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c112
*+ bl_0_112 br_0_112 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c112
*+ bl_0_112 br_0_112 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c112
*+ bl_0_112 br_0_112 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c112
*+ bl_0_112 br_0_112 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c112
*+ bl_0_112 br_0_112 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c112
*+ bl_0_112 br_0_112 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c112
*+ bl_0_112 br_0_112 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c112
*+ bl_0_112 br_0_112 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c112
*+ bl_0_112 br_0_112 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c112
*+ bl_0_112 br_0_112 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c112
*+ bl_0_112 br_0_112 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c112
*+ bl_0_112 br_0_112 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c112
*+ bl_0_112 br_0_112 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c112
*+ bl_0_112 br_0_112 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c112
*+ bl_0_112 br_0_112 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c112
*+ bl_0_112 br_0_112 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c112
*+ bl_0_112 br_0_112 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c112
*+ bl_0_112 br_0_112 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c112
*+ bl_0_112 br_0_112 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c112
*+ bl_0_112 br_0_112 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c112
*+ bl_0_112 br_0_112 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c112
*+ bl_0_112 br_0_112 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c112
*+ bl_0_112 br_0_112 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c112
*+ bl_0_112 br_0_112 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c112
*+ bl_0_112 br_0_112 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c112
*+ bl_0_112 br_0_112 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c112
*+ bl_0_112 br_0_112 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c112
*+ bl_0_112 br_0_112 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c112
*+ bl_0_112 br_0_112 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c112
*+ bl_0_112 br_0_112 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c112
*+ bl_0_112 br_0_112 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c112
*+ bl_0_112 br_0_112 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c112
*+ bl_0_112 br_0_112 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c112
*+ bl_0_112 br_0_112 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c112
*+ bl_0_112 br_0_112 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c112
*+ bl_0_112 br_0_112 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c112
*+ bl_0_112 br_0_112 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c112
*+ bl_0_112 br_0_112 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c112
*+ bl_0_112 br_0_112 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c112
*+ bl_0_112 br_0_112 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c112
*+ bl_0_112 br_0_112 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c112
*+ bl_0_112 br_0_112 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c112
*+ bl_0_112 br_0_112 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c112
*+ bl_0_112 br_0_112 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c112
*+ bl_0_112 br_0_112 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c112
*+ bl_0_112 br_0_112 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c112
*+ bl_0_112 br_0_112 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c112
*+ bl_0_112 br_0_112 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c112
*+ bl_0_112 br_0_112 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c112
*+ bl_0_112 br_0_112 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c112
*+ bl_0_112 br_0_112 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c112
*+ bl_0_112 br_0_112 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c112
*+ bl_0_112 br_0_112 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c112
*+ bl_0_112 br_0_112 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c112
*+ bl_0_112 br_0_112 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c112
*+ bl_0_112 br_0_112 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c112
*+ bl_0_112 br_0_112 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c112
*+ bl_0_112 br_0_112 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c112
*+ bl_0_112 br_0_112 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c112
*+ bl_0_112 br_0_112 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c112
*+ bl_0_112 br_0_112 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c112
*+ bl_0_112 br_0_112 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c112
*+ bl_0_112 br_0_112 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c112
*+ bl_0_112 br_0_112 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c112
*+ bl_0_112 br_0_112 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c112
*+ bl_0_112 br_0_112 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c112
*+ bl_0_112 br_0_112 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c112
*+ bl_0_112 br_0_112 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c112
*+ bl_0_112 br_0_112 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c112
*+ bl_0_112 br_0_112 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c112
*+ bl_0_112 br_0_112 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c112
*+ bl_0_112 br_0_112 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c112
+ bl_0_112 br_0_112 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c113
+ bl_0_113 br_0_113 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c113
*+ bl_0_113 br_0_113 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c113
*+ bl_0_113 br_0_113 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c113
*+ bl_0_113 br_0_113 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c113
*+ bl_0_113 br_0_113 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c113
*+ bl_0_113 br_0_113 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c113
*+ bl_0_113 br_0_113 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c113
*+ bl_0_113 br_0_113 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c113
*+ bl_0_113 br_0_113 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c113
*+ bl_0_113 br_0_113 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c113
*+ bl_0_113 br_0_113 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c113
*+ bl_0_113 br_0_113 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c113
*+ bl_0_113 br_0_113 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c113
*+ bl_0_113 br_0_113 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c113
*+ bl_0_113 br_0_113 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c113
*+ bl_0_113 br_0_113 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c113
*+ bl_0_113 br_0_113 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c113
*+ bl_0_113 br_0_113 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c113
*+ bl_0_113 br_0_113 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c113
*+ bl_0_113 br_0_113 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c113
*+ bl_0_113 br_0_113 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c113
*+ bl_0_113 br_0_113 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c113
*+ bl_0_113 br_0_113 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c113
*+ bl_0_113 br_0_113 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c113
*+ bl_0_113 br_0_113 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c113
*+ bl_0_113 br_0_113 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c113
*+ bl_0_113 br_0_113 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c113
*+ bl_0_113 br_0_113 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c113
*+ bl_0_113 br_0_113 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c113
*+ bl_0_113 br_0_113 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c113
*+ bl_0_113 br_0_113 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c113
*+ bl_0_113 br_0_113 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c113
*+ bl_0_113 br_0_113 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c113
*+ bl_0_113 br_0_113 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c113
*+ bl_0_113 br_0_113 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c113
*+ bl_0_113 br_0_113 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c113
*+ bl_0_113 br_0_113 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c113
*+ bl_0_113 br_0_113 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c113
*+ bl_0_113 br_0_113 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c113
*+ bl_0_113 br_0_113 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c113
*+ bl_0_113 br_0_113 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c113
*+ bl_0_113 br_0_113 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c113
*+ bl_0_113 br_0_113 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c113
*+ bl_0_113 br_0_113 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c113
*+ bl_0_113 br_0_113 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c113
*+ bl_0_113 br_0_113 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c113
*+ bl_0_113 br_0_113 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c113
*+ bl_0_113 br_0_113 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c113
*+ bl_0_113 br_0_113 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c113
*+ bl_0_113 br_0_113 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c113
*+ bl_0_113 br_0_113 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c113
*+ bl_0_113 br_0_113 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c113
*+ bl_0_113 br_0_113 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c113
*+ bl_0_113 br_0_113 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c113
*+ bl_0_113 br_0_113 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c113
*+ bl_0_113 br_0_113 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c113
*+ bl_0_113 br_0_113 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c113
*+ bl_0_113 br_0_113 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c113
*+ bl_0_113 br_0_113 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c113
*+ bl_0_113 br_0_113 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c113
*+ bl_0_113 br_0_113 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c113
*+ bl_0_113 br_0_113 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c113
*+ bl_0_113 br_0_113 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c113
*+ bl_0_113 br_0_113 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c113
*+ bl_0_113 br_0_113 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c113
*+ bl_0_113 br_0_113 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c113
*+ bl_0_113 br_0_113 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c113
*+ bl_0_113 br_0_113 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c113
*+ bl_0_113 br_0_113 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c113
*+ bl_0_113 br_0_113 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c113
*+ bl_0_113 br_0_113 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c113
*+ bl_0_113 br_0_113 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c113
*+ bl_0_113 br_0_113 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c113
*+ bl_0_113 br_0_113 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c113
*+ bl_0_113 br_0_113 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c113
*+ bl_0_113 br_0_113 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c113
*+ bl_0_113 br_0_113 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c113
*+ bl_0_113 br_0_113 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c113
*+ bl_0_113 br_0_113 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c113
*+ bl_0_113 br_0_113 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c113
*+ bl_0_113 br_0_113 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c113
*+ bl_0_113 br_0_113 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c113
*+ bl_0_113 br_0_113 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c113
*+ bl_0_113 br_0_113 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c113
*+ bl_0_113 br_0_113 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c113
*+ bl_0_113 br_0_113 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c113
*+ bl_0_113 br_0_113 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c113
*+ bl_0_113 br_0_113 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c113
*+ bl_0_113 br_0_113 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c113
*+ bl_0_113 br_0_113 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c113
*+ bl_0_113 br_0_113 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c113
*+ bl_0_113 br_0_113 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c113
*+ bl_0_113 br_0_113 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c113
*+ bl_0_113 br_0_113 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c113
*+ bl_0_113 br_0_113 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c113
*+ bl_0_113 br_0_113 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c113
*+ bl_0_113 br_0_113 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c113
*+ bl_0_113 br_0_113 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c113
*+ bl_0_113 br_0_113 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c113
*+ bl_0_113 br_0_113 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c113
*+ bl_0_113 br_0_113 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c113
*+ bl_0_113 br_0_113 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c113
*+ bl_0_113 br_0_113 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c113
*+ bl_0_113 br_0_113 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c113
*+ bl_0_113 br_0_113 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c113
*+ bl_0_113 br_0_113 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c113
*+ bl_0_113 br_0_113 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c113
*+ bl_0_113 br_0_113 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c113
*+ bl_0_113 br_0_113 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c113
*+ bl_0_113 br_0_113 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c113
*+ bl_0_113 br_0_113 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c113
*+ bl_0_113 br_0_113 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c113
*+ bl_0_113 br_0_113 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c113
*+ bl_0_113 br_0_113 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c113
*+ bl_0_113 br_0_113 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c113
*+ bl_0_113 br_0_113 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c113
*+ bl_0_113 br_0_113 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c113
*+ bl_0_113 br_0_113 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c113
*+ bl_0_113 br_0_113 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c113
*+ bl_0_113 br_0_113 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c113
*+ bl_0_113 br_0_113 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c113
*+ bl_0_113 br_0_113 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c113
*+ bl_0_113 br_0_113 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c113
*+ bl_0_113 br_0_113 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c113
*+ bl_0_113 br_0_113 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c113
*+ bl_0_113 br_0_113 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c113
*+ bl_0_113 br_0_113 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c113
+ bl_0_113 br_0_113 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c114
+ bl_0_114 br_0_114 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c114
*+ bl_0_114 br_0_114 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c114
*+ bl_0_114 br_0_114 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c114
*+ bl_0_114 br_0_114 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c114
*+ bl_0_114 br_0_114 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c114
*+ bl_0_114 br_0_114 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c114
*+ bl_0_114 br_0_114 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c114
*+ bl_0_114 br_0_114 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c114
*+ bl_0_114 br_0_114 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c114
*+ bl_0_114 br_0_114 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c114
*+ bl_0_114 br_0_114 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c114
*+ bl_0_114 br_0_114 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c114
*+ bl_0_114 br_0_114 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c114
*+ bl_0_114 br_0_114 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c114
*+ bl_0_114 br_0_114 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c114
*+ bl_0_114 br_0_114 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c114
*+ bl_0_114 br_0_114 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c114
*+ bl_0_114 br_0_114 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c114
*+ bl_0_114 br_0_114 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c114
*+ bl_0_114 br_0_114 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c114
*+ bl_0_114 br_0_114 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c114
*+ bl_0_114 br_0_114 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c114
*+ bl_0_114 br_0_114 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c114
*+ bl_0_114 br_0_114 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c114
*+ bl_0_114 br_0_114 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c114
*+ bl_0_114 br_0_114 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c114
*+ bl_0_114 br_0_114 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c114
*+ bl_0_114 br_0_114 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c114
*+ bl_0_114 br_0_114 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c114
*+ bl_0_114 br_0_114 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c114
*+ bl_0_114 br_0_114 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c114
*+ bl_0_114 br_0_114 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c114
*+ bl_0_114 br_0_114 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c114
*+ bl_0_114 br_0_114 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c114
*+ bl_0_114 br_0_114 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c114
*+ bl_0_114 br_0_114 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c114
*+ bl_0_114 br_0_114 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c114
*+ bl_0_114 br_0_114 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c114
*+ bl_0_114 br_0_114 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c114
*+ bl_0_114 br_0_114 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c114
*+ bl_0_114 br_0_114 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c114
*+ bl_0_114 br_0_114 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c114
*+ bl_0_114 br_0_114 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c114
*+ bl_0_114 br_0_114 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c114
*+ bl_0_114 br_0_114 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c114
*+ bl_0_114 br_0_114 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c114
*+ bl_0_114 br_0_114 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c114
*+ bl_0_114 br_0_114 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c114
*+ bl_0_114 br_0_114 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c114
*+ bl_0_114 br_0_114 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c114
*+ bl_0_114 br_0_114 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c114
*+ bl_0_114 br_0_114 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c114
*+ bl_0_114 br_0_114 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c114
*+ bl_0_114 br_0_114 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c114
*+ bl_0_114 br_0_114 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c114
*+ bl_0_114 br_0_114 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c114
*+ bl_0_114 br_0_114 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c114
*+ bl_0_114 br_0_114 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c114
*+ bl_0_114 br_0_114 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c114
*+ bl_0_114 br_0_114 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c114
*+ bl_0_114 br_0_114 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c114
*+ bl_0_114 br_0_114 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c114
*+ bl_0_114 br_0_114 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c114
*+ bl_0_114 br_0_114 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c114
*+ bl_0_114 br_0_114 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c114
*+ bl_0_114 br_0_114 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c114
*+ bl_0_114 br_0_114 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c114
*+ bl_0_114 br_0_114 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c114
*+ bl_0_114 br_0_114 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c114
*+ bl_0_114 br_0_114 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c114
*+ bl_0_114 br_0_114 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c114
*+ bl_0_114 br_0_114 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c114
*+ bl_0_114 br_0_114 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c114
*+ bl_0_114 br_0_114 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c114
*+ bl_0_114 br_0_114 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c114
*+ bl_0_114 br_0_114 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c114
*+ bl_0_114 br_0_114 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c114
*+ bl_0_114 br_0_114 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c114
*+ bl_0_114 br_0_114 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c114
*+ bl_0_114 br_0_114 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c114
*+ bl_0_114 br_0_114 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c114
*+ bl_0_114 br_0_114 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c114
*+ bl_0_114 br_0_114 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c114
*+ bl_0_114 br_0_114 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c114
*+ bl_0_114 br_0_114 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c114
*+ bl_0_114 br_0_114 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c114
*+ bl_0_114 br_0_114 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c114
*+ bl_0_114 br_0_114 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c114
*+ bl_0_114 br_0_114 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c114
*+ bl_0_114 br_0_114 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c114
*+ bl_0_114 br_0_114 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c114
*+ bl_0_114 br_0_114 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c114
*+ bl_0_114 br_0_114 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c114
*+ bl_0_114 br_0_114 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c114
*+ bl_0_114 br_0_114 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c114
*+ bl_0_114 br_0_114 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c114
*+ bl_0_114 br_0_114 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c114
*+ bl_0_114 br_0_114 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c114
*+ bl_0_114 br_0_114 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c114
*+ bl_0_114 br_0_114 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c114
*+ bl_0_114 br_0_114 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c114
*+ bl_0_114 br_0_114 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c114
*+ bl_0_114 br_0_114 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c114
*+ bl_0_114 br_0_114 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c114
*+ bl_0_114 br_0_114 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c114
*+ bl_0_114 br_0_114 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c114
*+ bl_0_114 br_0_114 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c114
*+ bl_0_114 br_0_114 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c114
*+ bl_0_114 br_0_114 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c114
*+ bl_0_114 br_0_114 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c114
*+ bl_0_114 br_0_114 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c114
*+ bl_0_114 br_0_114 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c114
*+ bl_0_114 br_0_114 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c114
*+ bl_0_114 br_0_114 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c114
*+ bl_0_114 br_0_114 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c114
*+ bl_0_114 br_0_114 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c114
*+ bl_0_114 br_0_114 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c114
*+ bl_0_114 br_0_114 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c114
*+ bl_0_114 br_0_114 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c114
*+ bl_0_114 br_0_114 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c114
*+ bl_0_114 br_0_114 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c114
*+ bl_0_114 br_0_114 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c114
*+ bl_0_114 br_0_114 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c114
*+ bl_0_114 br_0_114 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c114
*+ bl_0_114 br_0_114 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c114
*+ bl_0_114 br_0_114 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c114
*+ bl_0_114 br_0_114 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c114
+ bl_0_114 br_0_114 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c115
+ bl_0_115 br_0_115 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c115
*+ bl_0_115 br_0_115 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c115
*+ bl_0_115 br_0_115 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c115
*+ bl_0_115 br_0_115 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c115
*+ bl_0_115 br_0_115 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c115
*+ bl_0_115 br_0_115 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c115
*+ bl_0_115 br_0_115 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c115
*+ bl_0_115 br_0_115 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c115
*+ bl_0_115 br_0_115 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c115
*+ bl_0_115 br_0_115 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c115
*+ bl_0_115 br_0_115 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c115
*+ bl_0_115 br_0_115 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c115
*+ bl_0_115 br_0_115 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c115
*+ bl_0_115 br_0_115 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c115
*+ bl_0_115 br_0_115 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c115
*+ bl_0_115 br_0_115 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c115
*+ bl_0_115 br_0_115 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c115
*+ bl_0_115 br_0_115 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c115
*+ bl_0_115 br_0_115 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c115
*+ bl_0_115 br_0_115 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c115
*+ bl_0_115 br_0_115 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c115
*+ bl_0_115 br_0_115 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c115
*+ bl_0_115 br_0_115 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c115
*+ bl_0_115 br_0_115 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c115
*+ bl_0_115 br_0_115 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c115
*+ bl_0_115 br_0_115 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c115
*+ bl_0_115 br_0_115 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c115
*+ bl_0_115 br_0_115 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c115
*+ bl_0_115 br_0_115 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c115
*+ bl_0_115 br_0_115 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c115
*+ bl_0_115 br_0_115 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c115
*+ bl_0_115 br_0_115 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c115
*+ bl_0_115 br_0_115 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c115
*+ bl_0_115 br_0_115 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c115
*+ bl_0_115 br_0_115 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c115
*+ bl_0_115 br_0_115 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c115
*+ bl_0_115 br_0_115 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c115
*+ bl_0_115 br_0_115 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c115
*+ bl_0_115 br_0_115 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c115
*+ bl_0_115 br_0_115 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c115
*+ bl_0_115 br_0_115 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c115
*+ bl_0_115 br_0_115 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c115
*+ bl_0_115 br_0_115 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c115
*+ bl_0_115 br_0_115 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c115
*+ bl_0_115 br_0_115 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c115
*+ bl_0_115 br_0_115 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c115
*+ bl_0_115 br_0_115 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c115
*+ bl_0_115 br_0_115 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c115
*+ bl_0_115 br_0_115 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c115
*+ bl_0_115 br_0_115 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c115
*+ bl_0_115 br_0_115 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c115
*+ bl_0_115 br_0_115 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c115
*+ bl_0_115 br_0_115 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c115
*+ bl_0_115 br_0_115 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c115
*+ bl_0_115 br_0_115 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c115
*+ bl_0_115 br_0_115 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c115
*+ bl_0_115 br_0_115 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c115
*+ bl_0_115 br_0_115 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c115
*+ bl_0_115 br_0_115 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c115
*+ bl_0_115 br_0_115 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c115
*+ bl_0_115 br_0_115 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c115
*+ bl_0_115 br_0_115 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c115
*+ bl_0_115 br_0_115 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c115
*+ bl_0_115 br_0_115 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c115
*+ bl_0_115 br_0_115 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c115
*+ bl_0_115 br_0_115 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c115
*+ bl_0_115 br_0_115 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c115
*+ bl_0_115 br_0_115 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c115
*+ bl_0_115 br_0_115 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c115
*+ bl_0_115 br_0_115 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c115
*+ bl_0_115 br_0_115 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c115
*+ bl_0_115 br_0_115 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c115
*+ bl_0_115 br_0_115 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c115
*+ bl_0_115 br_0_115 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c115
*+ bl_0_115 br_0_115 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c115
*+ bl_0_115 br_0_115 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c115
*+ bl_0_115 br_0_115 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c115
*+ bl_0_115 br_0_115 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c115
*+ bl_0_115 br_0_115 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c115
*+ bl_0_115 br_0_115 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c115
*+ bl_0_115 br_0_115 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c115
*+ bl_0_115 br_0_115 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c115
*+ bl_0_115 br_0_115 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c115
*+ bl_0_115 br_0_115 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c115
*+ bl_0_115 br_0_115 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c115
*+ bl_0_115 br_0_115 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c115
*+ bl_0_115 br_0_115 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c115
*+ bl_0_115 br_0_115 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c115
*+ bl_0_115 br_0_115 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c115
*+ bl_0_115 br_0_115 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c115
*+ bl_0_115 br_0_115 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c115
*+ bl_0_115 br_0_115 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c115
*+ bl_0_115 br_0_115 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c115
*+ bl_0_115 br_0_115 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c115
*+ bl_0_115 br_0_115 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c115
*+ bl_0_115 br_0_115 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c115
*+ bl_0_115 br_0_115 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c115
*+ bl_0_115 br_0_115 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c115
*+ bl_0_115 br_0_115 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c115
*+ bl_0_115 br_0_115 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c115
*+ bl_0_115 br_0_115 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c115
*+ bl_0_115 br_0_115 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c115
*+ bl_0_115 br_0_115 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c115
*+ bl_0_115 br_0_115 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c115
*+ bl_0_115 br_0_115 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c115
*+ bl_0_115 br_0_115 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c115
*+ bl_0_115 br_0_115 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c115
*+ bl_0_115 br_0_115 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c115
*+ bl_0_115 br_0_115 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c115
*+ bl_0_115 br_0_115 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c115
*+ bl_0_115 br_0_115 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c115
*+ bl_0_115 br_0_115 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c115
*+ bl_0_115 br_0_115 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c115
*+ bl_0_115 br_0_115 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c115
*+ bl_0_115 br_0_115 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c115
*+ bl_0_115 br_0_115 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c115
*+ bl_0_115 br_0_115 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c115
*+ bl_0_115 br_0_115 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c115
*+ bl_0_115 br_0_115 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c115
*+ bl_0_115 br_0_115 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c115
*+ bl_0_115 br_0_115 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c115
*+ bl_0_115 br_0_115 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c115
*+ bl_0_115 br_0_115 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c115
*+ bl_0_115 br_0_115 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c115
*+ bl_0_115 br_0_115 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c115
*+ bl_0_115 br_0_115 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c115
*+ bl_0_115 br_0_115 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c115
+ bl_0_115 br_0_115 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c116
+ bl_0_116 br_0_116 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c116
*+ bl_0_116 br_0_116 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c116
*+ bl_0_116 br_0_116 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c116
*+ bl_0_116 br_0_116 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c116
*+ bl_0_116 br_0_116 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c116
*+ bl_0_116 br_0_116 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c116
*+ bl_0_116 br_0_116 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c116
*+ bl_0_116 br_0_116 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c116
*+ bl_0_116 br_0_116 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c116
*+ bl_0_116 br_0_116 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c116
*+ bl_0_116 br_0_116 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c116
*+ bl_0_116 br_0_116 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c116
*+ bl_0_116 br_0_116 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c116
*+ bl_0_116 br_0_116 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c116
*+ bl_0_116 br_0_116 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c116
*+ bl_0_116 br_0_116 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c116
*+ bl_0_116 br_0_116 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c116
*+ bl_0_116 br_0_116 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c116
*+ bl_0_116 br_0_116 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c116
*+ bl_0_116 br_0_116 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c116
*+ bl_0_116 br_0_116 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c116
*+ bl_0_116 br_0_116 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c116
*+ bl_0_116 br_0_116 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c116
*+ bl_0_116 br_0_116 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c116
*+ bl_0_116 br_0_116 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c116
*+ bl_0_116 br_0_116 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c116
*+ bl_0_116 br_0_116 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c116
*+ bl_0_116 br_0_116 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c116
*+ bl_0_116 br_0_116 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c116
*+ bl_0_116 br_0_116 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c116
*+ bl_0_116 br_0_116 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c116
*+ bl_0_116 br_0_116 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c116
*+ bl_0_116 br_0_116 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c116
*+ bl_0_116 br_0_116 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c116
*+ bl_0_116 br_0_116 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c116
*+ bl_0_116 br_0_116 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c116
*+ bl_0_116 br_0_116 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c116
*+ bl_0_116 br_0_116 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c116
*+ bl_0_116 br_0_116 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c116
*+ bl_0_116 br_0_116 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c116
*+ bl_0_116 br_0_116 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c116
*+ bl_0_116 br_0_116 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c116
*+ bl_0_116 br_0_116 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c116
*+ bl_0_116 br_0_116 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c116
*+ bl_0_116 br_0_116 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c116
*+ bl_0_116 br_0_116 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c116
*+ bl_0_116 br_0_116 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c116
*+ bl_0_116 br_0_116 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c116
*+ bl_0_116 br_0_116 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c116
*+ bl_0_116 br_0_116 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c116
*+ bl_0_116 br_0_116 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c116
*+ bl_0_116 br_0_116 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c116
*+ bl_0_116 br_0_116 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c116
*+ bl_0_116 br_0_116 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c116
*+ bl_0_116 br_0_116 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c116
*+ bl_0_116 br_0_116 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c116
*+ bl_0_116 br_0_116 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c116
*+ bl_0_116 br_0_116 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c116
*+ bl_0_116 br_0_116 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c116
*+ bl_0_116 br_0_116 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c116
*+ bl_0_116 br_0_116 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c116
*+ bl_0_116 br_0_116 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c116
*+ bl_0_116 br_0_116 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c116
*+ bl_0_116 br_0_116 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c116
*+ bl_0_116 br_0_116 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c116
*+ bl_0_116 br_0_116 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c116
*+ bl_0_116 br_0_116 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c116
*+ bl_0_116 br_0_116 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c116
*+ bl_0_116 br_0_116 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c116
*+ bl_0_116 br_0_116 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c116
*+ bl_0_116 br_0_116 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c116
*+ bl_0_116 br_0_116 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c116
*+ bl_0_116 br_0_116 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c116
*+ bl_0_116 br_0_116 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c116
*+ bl_0_116 br_0_116 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c116
*+ bl_0_116 br_0_116 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c116
*+ bl_0_116 br_0_116 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c116
*+ bl_0_116 br_0_116 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c116
*+ bl_0_116 br_0_116 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c116
*+ bl_0_116 br_0_116 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c116
*+ bl_0_116 br_0_116 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c116
*+ bl_0_116 br_0_116 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c116
*+ bl_0_116 br_0_116 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c116
*+ bl_0_116 br_0_116 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c116
*+ bl_0_116 br_0_116 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c116
*+ bl_0_116 br_0_116 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c116
*+ bl_0_116 br_0_116 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c116
*+ bl_0_116 br_0_116 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c116
*+ bl_0_116 br_0_116 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c116
*+ bl_0_116 br_0_116 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c116
*+ bl_0_116 br_0_116 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c116
*+ bl_0_116 br_0_116 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c116
*+ bl_0_116 br_0_116 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c116
*+ bl_0_116 br_0_116 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c116
*+ bl_0_116 br_0_116 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c116
*+ bl_0_116 br_0_116 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c116
*+ bl_0_116 br_0_116 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c116
*+ bl_0_116 br_0_116 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c116
*+ bl_0_116 br_0_116 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c116
*+ bl_0_116 br_0_116 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c116
*+ bl_0_116 br_0_116 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c116
*+ bl_0_116 br_0_116 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c116
*+ bl_0_116 br_0_116 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c116
*+ bl_0_116 br_0_116 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c116
*+ bl_0_116 br_0_116 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c116
*+ bl_0_116 br_0_116 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c116
*+ bl_0_116 br_0_116 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c116
*+ bl_0_116 br_0_116 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c116
*+ bl_0_116 br_0_116 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c116
*+ bl_0_116 br_0_116 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c116
*+ bl_0_116 br_0_116 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c116
*+ bl_0_116 br_0_116 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c116
*+ bl_0_116 br_0_116 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c116
*+ bl_0_116 br_0_116 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c116
*+ bl_0_116 br_0_116 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c116
*+ bl_0_116 br_0_116 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c116
*+ bl_0_116 br_0_116 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c116
*+ bl_0_116 br_0_116 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c116
*+ bl_0_116 br_0_116 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c116
*+ bl_0_116 br_0_116 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c116
*+ bl_0_116 br_0_116 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c116
*+ bl_0_116 br_0_116 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c116
*+ bl_0_116 br_0_116 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c116
*+ bl_0_116 br_0_116 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c116
*+ bl_0_116 br_0_116 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c116
*+ bl_0_116 br_0_116 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c116
*+ bl_0_116 br_0_116 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c116
+ bl_0_116 br_0_116 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c117
+ bl_0_117 br_0_117 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c117
*+ bl_0_117 br_0_117 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c117
*+ bl_0_117 br_0_117 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c117
*+ bl_0_117 br_0_117 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c117
*+ bl_0_117 br_0_117 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c117
*+ bl_0_117 br_0_117 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c117
*+ bl_0_117 br_0_117 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c117
*+ bl_0_117 br_0_117 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c117
*+ bl_0_117 br_0_117 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c117
*+ bl_0_117 br_0_117 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c117
*+ bl_0_117 br_0_117 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c117
*+ bl_0_117 br_0_117 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c117
*+ bl_0_117 br_0_117 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c117
*+ bl_0_117 br_0_117 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c117
*+ bl_0_117 br_0_117 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c117
*+ bl_0_117 br_0_117 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c117
*+ bl_0_117 br_0_117 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c117
*+ bl_0_117 br_0_117 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c117
*+ bl_0_117 br_0_117 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c117
*+ bl_0_117 br_0_117 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c117
*+ bl_0_117 br_0_117 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c117
*+ bl_0_117 br_0_117 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c117
*+ bl_0_117 br_0_117 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c117
*+ bl_0_117 br_0_117 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c117
*+ bl_0_117 br_0_117 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c117
*+ bl_0_117 br_0_117 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c117
*+ bl_0_117 br_0_117 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c117
*+ bl_0_117 br_0_117 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c117
*+ bl_0_117 br_0_117 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c117
*+ bl_0_117 br_0_117 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c117
*+ bl_0_117 br_0_117 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c117
*+ bl_0_117 br_0_117 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c117
*+ bl_0_117 br_0_117 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c117
*+ bl_0_117 br_0_117 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c117
*+ bl_0_117 br_0_117 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c117
*+ bl_0_117 br_0_117 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c117
*+ bl_0_117 br_0_117 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c117
*+ bl_0_117 br_0_117 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c117
*+ bl_0_117 br_0_117 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c117
*+ bl_0_117 br_0_117 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c117
*+ bl_0_117 br_0_117 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c117
*+ bl_0_117 br_0_117 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c117
*+ bl_0_117 br_0_117 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c117
*+ bl_0_117 br_0_117 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c117
*+ bl_0_117 br_0_117 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c117
*+ bl_0_117 br_0_117 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c117
*+ bl_0_117 br_0_117 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c117
*+ bl_0_117 br_0_117 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c117
*+ bl_0_117 br_0_117 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c117
*+ bl_0_117 br_0_117 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c117
*+ bl_0_117 br_0_117 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c117
*+ bl_0_117 br_0_117 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c117
*+ bl_0_117 br_0_117 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c117
*+ bl_0_117 br_0_117 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c117
*+ bl_0_117 br_0_117 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c117
*+ bl_0_117 br_0_117 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c117
*+ bl_0_117 br_0_117 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c117
*+ bl_0_117 br_0_117 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c117
*+ bl_0_117 br_0_117 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c117
*+ bl_0_117 br_0_117 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c117
*+ bl_0_117 br_0_117 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c117
*+ bl_0_117 br_0_117 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c117
*+ bl_0_117 br_0_117 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c117
*+ bl_0_117 br_0_117 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c117
*+ bl_0_117 br_0_117 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c117
*+ bl_0_117 br_0_117 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c117
*+ bl_0_117 br_0_117 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c117
*+ bl_0_117 br_0_117 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c117
*+ bl_0_117 br_0_117 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c117
*+ bl_0_117 br_0_117 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c117
*+ bl_0_117 br_0_117 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c117
*+ bl_0_117 br_0_117 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c117
*+ bl_0_117 br_0_117 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c117
*+ bl_0_117 br_0_117 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c117
*+ bl_0_117 br_0_117 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c117
*+ bl_0_117 br_0_117 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c117
*+ bl_0_117 br_0_117 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c117
*+ bl_0_117 br_0_117 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c117
*+ bl_0_117 br_0_117 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c117
*+ bl_0_117 br_0_117 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c117
*+ bl_0_117 br_0_117 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c117
*+ bl_0_117 br_0_117 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c117
*+ bl_0_117 br_0_117 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c117
*+ bl_0_117 br_0_117 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c117
*+ bl_0_117 br_0_117 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c117
*+ bl_0_117 br_0_117 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c117
*+ bl_0_117 br_0_117 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c117
*+ bl_0_117 br_0_117 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c117
*+ bl_0_117 br_0_117 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c117
*+ bl_0_117 br_0_117 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c117
*+ bl_0_117 br_0_117 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c117
*+ bl_0_117 br_0_117 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c117
*+ bl_0_117 br_0_117 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c117
*+ bl_0_117 br_0_117 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c117
*+ bl_0_117 br_0_117 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c117
*+ bl_0_117 br_0_117 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c117
*+ bl_0_117 br_0_117 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c117
*+ bl_0_117 br_0_117 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c117
*+ bl_0_117 br_0_117 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c117
*+ bl_0_117 br_0_117 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c117
*+ bl_0_117 br_0_117 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c117
*+ bl_0_117 br_0_117 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c117
*+ bl_0_117 br_0_117 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c117
*+ bl_0_117 br_0_117 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c117
*+ bl_0_117 br_0_117 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c117
*+ bl_0_117 br_0_117 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c117
*+ bl_0_117 br_0_117 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c117
*+ bl_0_117 br_0_117 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c117
*+ bl_0_117 br_0_117 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c117
*+ bl_0_117 br_0_117 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c117
*+ bl_0_117 br_0_117 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c117
*+ bl_0_117 br_0_117 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c117
*+ bl_0_117 br_0_117 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c117
*+ bl_0_117 br_0_117 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c117
*+ bl_0_117 br_0_117 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c117
*+ bl_0_117 br_0_117 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c117
*+ bl_0_117 br_0_117 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c117
*+ bl_0_117 br_0_117 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c117
*+ bl_0_117 br_0_117 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c117
*+ bl_0_117 br_0_117 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c117
*+ bl_0_117 br_0_117 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c117
*+ bl_0_117 br_0_117 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c117
*+ bl_0_117 br_0_117 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c117
*+ bl_0_117 br_0_117 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c117
*+ bl_0_117 br_0_117 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c117
*+ bl_0_117 br_0_117 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c117
*+ bl_0_117 br_0_117 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c117
+ bl_0_117 br_0_117 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c118
+ bl_0_118 br_0_118 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c118
*+ bl_0_118 br_0_118 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c118
*+ bl_0_118 br_0_118 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c118
*+ bl_0_118 br_0_118 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c118
*+ bl_0_118 br_0_118 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c118
*+ bl_0_118 br_0_118 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c118
*+ bl_0_118 br_0_118 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c118
*+ bl_0_118 br_0_118 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c118
*+ bl_0_118 br_0_118 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c118
*+ bl_0_118 br_0_118 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c118
*+ bl_0_118 br_0_118 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c118
*+ bl_0_118 br_0_118 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c118
*+ bl_0_118 br_0_118 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c118
*+ bl_0_118 br_0_118 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c118
*+ bl_0_118 br_0_118 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c118
*+ bl_0_118 br_0_118 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c118
*+ bl_0_118 br_0_118 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c118
*+ bl_0_118 br_0_118 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c118
*+ bl_0_118 br_0_118 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c118
*+ bl_0_118 br_0_118 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c118
*+ bl_0_118 br_0_118 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c118
*+ bl_0_118 br_0_118 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c118
*+ bl_0_118 br_0_118 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c118
*+ bl_0_118 br_0_118 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c118
*+ bl_0_118 br_0_118 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c118
*+ bl_0_118 br_0_118 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c118
*+ bl_0_118 br_0_118 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c118
*+ bl_0_118 br_0_118 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c118
*+ bl_0_118 br_0_118 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c118
*+ bl_0_118 br_0_118 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c118
*+ bl_0_118 br_0_118 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c118
*+ bl_0_118 br_0_118 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c118
*+ bl_0_118 br_0_118 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c118
*+ bl_0_118 br_0_118 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c118
*+ bl_0_118 br_0_118 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c118
*+ bl_0_118 br_0_118 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c118
*+ bl_0_118 br_0_118 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c118
*+ bl_0_118 br_0_118 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c118
*+ bl_0_118 br_0_118 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c118
*+ bl_0_118 br_0_118 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c118
*+ bl_0_118 br_0_118 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c118
*+ bl_0_118 br_0_118 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c118
*+ bl_0_118 br_0_118 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c118
*+ bl_0_118 br_0_118 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c118
*+ bl_0_118 br_0_118 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c118
*+ bl_0_118 br_0_118 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c118
*+ bl_0_118 br_0_118 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c118
*+ bl_0_118 br_0_118 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c118
*+ bl_0_118 br_0_118 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c118
*+ bl_0_118 br_0_118 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c118
*+ bl_0_118 br_0_118 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c118
*+ bl_0_118 br_0_118 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c118
*+ bl_0_118 br_0_118 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c118
*+ bl_0_118 br_0_118 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c118
*+ bl_0_118 br_0_118 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c118
*+ bl_0_118 br_0_118 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c118
*+ bl_0_118 br_0_118 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c118
*+ bl_0_118 br_0_118 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c118
*+ bl_0_118 br_0_118 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c118
*+ bl_0_118 br_0_118 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c118
*+ bl_0_118 br_0_118 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c118
*+ bl_0_118 br_0_118 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c118
*+ bl_0_118 br_0_118 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c118
*+ bl_0_118 br_0_118 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c118
*+ bl_0_118 br_0_118 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c118
*+ bl_0_118 br_0_118 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c118
*+ bl_0_118 br_0_118 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c118
*+ bl_0_118 br_0_118 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c118
*+ bl_0_118 br_0_118 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c118
*+ bl_0_118 br_0_118 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c118
*+ bl_0_118 br_0_118 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c118
*+ bl_0_118 br_0_118 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c118
*+ bl_0_118 br_0_118 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c118
*+ bl_0_118 br_0_118 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c118
*+ bl_0_118 br_0_118 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c118
*+ bl_0_118 br_0_118 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c118
*+ bl_0_118 br_0_118 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c118
*+ bl_0_118 br_0_118 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c118
*+ bl_0_118 br_0_118 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c118
*+ bl_0_118 br_0_118 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c118
*+ bl_0_118 br_0_118 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c118
*+ bl_0_118 br_0_118 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c118
*+ bl_0_118 br_0_118 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c118
*+ bl_0_118 br_0_118 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c118
*+ bl_0_118 br_0_118 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c118
*+ bl_0_118 br_0_118 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c118
*+ bl_0_118 br_0_118 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c118
*+ bl_0_118 br_0_118 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c118
*+ bl_0_118 br_0_118 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c118
*+ bl_0_118 br_0_118 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c118
*+ bl_0_118 br_0_118 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c118
*+ bl_0_118 br_0_118 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c118
*+ bl_0_118 br_0_118 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c118
*+ bl_0_118 br_0_118 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c118
*+ bl_0_118 br_0_118 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c118
*+ bl_0_118 br_0_118 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c118
*+ bl_0_118 br_0_118 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c118
*+ bl_0_118 br_0_118 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c118
*+ bl_0_118 br_0_118 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c118
*+ bl_0_118 br_0_118 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c118
*+ bl_0_118 br_0_118 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c118
*+ bl_0_118 br_0_118 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c118
*+ bl_0_118 br_0_118 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c118
*+ bl_0_118 br_0_118 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c118
*+ bl_0_118 br_0_118 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c118
*+ bl_0_118 br_0_118 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c118
*+ bl_0_118 br_0_118 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c118
*+ bl_0_118 br_0_118 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c118
*+ bl_0_118 br_0_118 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c118
*+ bl_0_118 br_0_118 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c118
*+ bl_0_118 br_0_118 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c118
*+ bl_0_118 br_0_118 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c118
*+ bl_0_118 br_0_118 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c118
*+ bl_0_118 br_0_118 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c118
*+ bl_0_118 br_0_118 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c118
*+ bl_0_118 br_0_118 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c118
*+ bl_0_118 br_0_118 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c118
*+ bl_0_118 br_0_118 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c118
*+ bl_0_118 br_0_118 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c118
*+ bl_0_118 br_0_118 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c118
*+ bl_0_118 br_0_118 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c118
*+ bl_0_118 br_0_118 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c118
*+ bl_0_118 br_0_118 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c118
*+ bl_0_118 br_0_118 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c118
*+ bl_0_118 br_0_118 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c118
*+ bl_0_118 br_0_118 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c118
*+ bl_0_118 br_0_118 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c118
+ bl_0_118 br_0_118 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c119
+ bl_0_119 br_0_119 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c119
*+ bl_0_119 br_0_119 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c119
*+ bl_0_119 br_0_119 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c119
*+ bl_0_119 br_0_119 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c119
*+ bl_0_119 br_0_119 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c119
*+ bl_0_119 br_0_119 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c119
*+ bl_0_119 br_0_119 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c119
*+ bl_0_119 br_0_119 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c119
*+ bl_0_119 br_0_119 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c119
*+ bl_0_119 br_0_119 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c119
*+ bl_0_119 br_0_119 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c119
*+ bl_0_119 br_0_119 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c119
*+ bl_0_119 br_0_119 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c119
*+ bl_0_119 br_0_119 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c119
*+ bl_0_119 br_0_119 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c119
*+ bl_0_119 br_0_119 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c119
*+ bl_0_119 br_0_119 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c119
*+ bl_0_119 br_0_119 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c119
*+ bl_0_119 br_0_119 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c119
*+ bl_0_119 br_0_119 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c119
*+ bl_0_119 br_0_119 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c119
*+ bl_0_119 br_0_119 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c119
*+ bl_0_119 br_0_119 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c119
*+ bl_0_119 br_0_119 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c119
*+ bl_0_119 br_0_119 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c119
*+ bl_0_119 br_0_119 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c119
*+ bl_0_119 br_0_119 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c119
*+ bl_0_119 br_0_119 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c119
*+ bl_0_119 br_0_119 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c119
*+ bl_0_119 br_0_119 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c119
*+ bl_0_119 br_0_119 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c119
*+ bl_0_119 br_0_119 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c119
*+ bl_0_119 br_0_119 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c119
*+ bl_0_119 br_0_119 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c119
*+ bl_0_119 br_0_119 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c119
*+ bl_0_119 br_0_119 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c119
*+ bl_0_119 br_0_119 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c119
*+ bl_0_119 br_0_119 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c119
*+ bl_0_119 br_0_119 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c119
*+ bl_0_119 br_0_119 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c119
*+ bl_0_119 br_0_119 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c119
*+ bl_0_119 br_0_119 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c119
*+ bl_0_119 br_0_119 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c119
*+ bl_0_119 br_0_119 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c119
*+ bl_0_119 br_0_119 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c119
*+ bl_0_119 br_0_119 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c119
*+ bl_0_119 br_0_119 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c119
*+ bl_0_119 br_0_119 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c119
*+ bl_0_119 br_0_119 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c119
*+ bl_0_119 br_0_119 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c119
*+ bl_0_119 br_0_119 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c119
*+ bl_0_119 br_0_119 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c119
*+ bl_0_119 br_0_119 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c119
*+ bl_0_119 br_0_119 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c119
*+ bl_0_119 br_0_119 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c119
*+ bl_0_119 br_0_119 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c119
*+ bl_0_119 br_0_119 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c119
*+ bl_0_119 br_0_119 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c119
*+ bl_0_119 br_0_119 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c119
*+ bl_0_119 br_0_119 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c119
*+ bl_0_119 br_0_119 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c119
*+ bl_0_119 br_0_119 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c119
*+ bl_0_119 br_0_119 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c119
*+ bl_0_119 br_0_119 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c119
*+ bl_0_119 br_0_119 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c119
*+ bl_0_119 br_0_119 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c119
*+ bl_0_119 br_0_119 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c119
*+ bl_0_119 br_0_119 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c119
*+ bl_0_119 br_0_119 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c119
*+ bl_0_119 br_0_119 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c119
*+ bl_0_119 br_0_119 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c119
*+ bl_0_119 br_0_119 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c119
*+ bl_0_119 br_0_119 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c119
*+ bl_0_119 br_0_119 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c119
*+ bl_0_119 br_0_119 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c119
*+ bl_0_119 br_0_119 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c119
*+ bl_0_119 br_0_119 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c119
*+ bl_0_119 br_0_119 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c119
*+ bl_0_119 br_0_119 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c119
*+ bl_0_119 br_0_119 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c119
*+ bl_0_119 br_0_119 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c119
*+ bl_0_119 br_0_119 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c119
*+ bl_0_119 br_0_119 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c119
*+ bl_0_119 br_0_119 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c119
*+ bl_0_119 br_0_119 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c119
*+ bl_0_119 br_0_119 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c119
*+ bl_0_119 br_0_119 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c119
*+ bl_0_119 br_0_119 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c119
*+ bl_0_119 br_0_119 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c119
*+ bl_0_119 br_0_119 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c119
*+ bl_0_119 br_0_119 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c119
*+ bl_0_119 br_0_119 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c119
*+ bl_0_119 br_0_119 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c119
*+ bl_0_119 br_0_119 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c119
*+ bl_0_119 br_0_119 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c119
*+ bl_0_119 br_0_119 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c119
*+ bl_0_119 br_0_119 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c119
*+ bl_0_119 br_0_119 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c119
*+ bl_0_119 br_0_119 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c119
*+ bl_0_119 br_0_119 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c119
*+ bl_0_119 br_0_119 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c119
*+ bl_0_119 br_0_119 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c119
*+ bl_0_119 br_0_119 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c119
*+ bl_0_119 br_0_119 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c119
*+ bl_0_119 br_0_119 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c119
*+ bl_0_119 br_0_119 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c119
*+ bl_0_119 br_0_119 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c119
*+ bl_0_119 br_0_119 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c119
*+ bl_0_119 br_0_119 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c119
*+ bl_0_119 br_0_119 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c119
*+ bl_0_119 br_0_119 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c119
*+ bl_0_119 br_0_119 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c119
*+ bl_0_119 br_0_119 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c119
*+ bl_0_119 br_0_119 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c119
*+ bl_0_119 br_0_119 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c119
*+ bl_0_119 br_0_119 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c119
*+ bl_0_119 br_0_119 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c119
*+ bl_0_119 br_0_119 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c119
*+ bl_0_119 br_0_119 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c119
*+ bl_0_119 br_0_119 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c119
*+ bl_0_119 br_0_119 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c119
*+ bl_0_119 br_0_119 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c119
*+ bl_0_119 br_0_119 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c119
*+ bl_0_119 br_0_119 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c119
*+ bl_0_119 br_0_119 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c119
*+ bl_0_119 br_0_119 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c119
*+ bl_0_119 br_0_119 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c119
+ bl_0_119 br_0_119 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c120
+ bl_0_120 br_0_120 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c120
*+ bl_0_120 br_0_120 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c120
*+ bl_0_120 br_0_120 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c120
*+ bl_0_120 br_0_120 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c120
*+ bl_0_120 br_0_120 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c120
*+ bl_0_120 br_0_120 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c120
*+ bl_0_120 br_0_120 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c120
*+ bl_0_120 br_0_120 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c120
*+ bl_0_120 br_0_120 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c120
*+ bl_0_120 br_0_120 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c120
*+ bl_0_120 br_0_120 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c120
*+ bl_0_120 br_0_120 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c120
*+ bl_0_120 br_0_120 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c120
*+ bl_0_120 br_0_120 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c120
*+ bl_0_120 br_0_120 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c120
*+ bl_0_120 br_0_120 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c120
*+ bl_0_120 br_0_120 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c120
*+ bl_0_120 br_0_120 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c120
*+ bl_0_120 br_0_120 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c120
*+ bl_0_120 br_0_120 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c120
*+ bl_0_120 br_0_120 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c120
*+ bl_0_120 br_0_120 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c120
*+ bl_0_120 br_0_120 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c120
*+ bl_0_120 br_0_120 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c120
*+ bl_0_120 br_0_120 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c120
*+ bl_0_120 br_0_120 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c120
*+ bl_0_120 br_0_120 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c120
*+ bl_0_120 br_0_120 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c120
*+ bl_0_120 br_0_120 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c120
*+ bl_0_120 br_0_120 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c120
*+ bl_0_120 br_0_120 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c120
*+ bl_0_120 br_0_120 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c120
*+ bl_0_120 br_0_120 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c120
*+ bl_0_120 br_0_120 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c120
*+ bl_0_120 br_0_120 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c120
*+ bl_0_120 br_0_120 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c120
*+ bl_0_120 br_0_120 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c120
*+ bl_0_120 br_0_120 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c120
*+ bl_0_120 br_0_120 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c120
*+ bl_0_120 br_0_120 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c120
*+ bl_0_120 br_0_120 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c120
*+ bl_0_120 br_0_120 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c120
*+ bl_0_120 br_0_120 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c120
*+ bl_0_120 br_0_120 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c120
*+ bl_0_120 br_0_120 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c120
*+ bl_0_120 br_0_120 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c120
*+ bl_0_120 br_0_120 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c120
*+ bl_0_120 br_0_120 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c120
*+ bl_0_120 br_0_120 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c120
*+ bl_0_120 br_0_120 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c120
*+ bl_0_120 br_0_120 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c120
*+ bl_0_120 br_0_120 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c120
*+ bl_0_120 br_0_120 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c120
*+ bl_0_120 br_0_120 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c120
*+ bl_0_120 br_0_120 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c120
*+ bl_0_120 br_0_120 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c120
*+ bl_0_120 br_0_120 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c120
*+ bl_0_120 br_0_120 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c120
*+ bl_0_120 br_0_120 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c120
*+ bl_0_120 br_0_120 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c120
*+ bl_0_120 br_0_120 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c120
*+ bl_0_120 br_0_120 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c120
*+ bl_0_120 br_0_120 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c120
*+ bl_0_120 br_0_120 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c120
*+ bl_0_120 br_0_120 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c120
*+ bl_0_120 br_0_120 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c120
*+ bl_0_120 br_0_120 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c120
*+ bl_0_120 br_0_120 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c120
*+ bl_0_120 br_0_120 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c120
*+ bl_0_120 br_0_120 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c120
*+ bl_0_120 br_0_120 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c120
*+ bl_0_120 br_0_120 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c120
*+ bl_0_120 br_0_120 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c120
*+ bl_0_120 br_0_120 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c120
*+ bl_0_120 br_0_120 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c120
*+ bl_0_120 br_0_120 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c120
*+ bl_0_120 br_0_120 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c120
*+ bl_0_120 br_0_120 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c120
*+ bl_0_120 br_0_120 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c120
*+ bl_0_120 br_0_120 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c120
*+ bl_0_120 br_0_120 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c120
*+ bl_0_120 br_0_120 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c120
*+ bl_0_120 br_0_120 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c120
*+ bl_0_120 br_0_120 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c120
*+ bl_0_120 br_0_120 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c120
*+ bl_0_120 br_0_120 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c120
*+ bl_0_120 br_0_120 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c120
*+ bl_0_120 br_0_120 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c120
*+ bl_0_120 br_0_120 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c120
*+ bl_0_120 br_0_120 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c120
*+ bl_0_120 br_0_120 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c120
*+ bl_0_120 br_0_120 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c120
*+ bl_0_120 br_0_120 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c120
*+ bl_0_120 br_0_120 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c120
*+ bl_0_120 br_0_120 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c120
*+ bl_0_120 br_0_120 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c120
*+ bl_0_120 br_0_120 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c120
*+ bl_0_120 br_0_120 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c120
*+ bl_0_120 br_0_120 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c120
*+ bl_0_120 br_0_120 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c120
*+ bl_0_120 br_0_120 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c120
*+ bl_0_120 br_0_120 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c120
*+ bl_0_120 br_0_120 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c120
*+ bl_0_120 br_0_120 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c120
*+ bl_0_120 br_0_120 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c120
*+ bl_0_120 br_0_120 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c120
*+ bl_0_120 br_0_120 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c120
*+ bl_0_120 br_0_120 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c120
*+ bl_0_120 br_0_120 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c120
*+ bl_0_120 br_0_120 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c120
*+ bl_0_120 br_0_120 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c120
*+ bl_0_120 br_0_120 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c120
*+ bl_0_120 br_0_120 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c120
*+ bl_0_120 br_0_120 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c120
*+ bl_0_120 br_0_120 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c120
*+ bl_0_120 br_0_120 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c120
*+ bl_0_120 br_0_120 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c120
*+ bl_0_120 br_0_120 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c120
*+ bl_0_120 br_0_120 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c120
*+ bl_0_120 br_0_120 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c120
*+ bl_0_120 br_0_120 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c120
*+ bl_0_120 br_0_120 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c120
*+ bl_0_120 br_0_120 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c120
*+ bl_0_120 br_0_120 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c120
*+ bl_0_120 br_0_120 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c120
*+ bl_0_120 br_0_120 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c120
*+ bl_0_120 br_0_120 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c120
+ bl_0_120 br_0_120 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c121
+ bl_0_121 br_0_121 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c121
*+ bl_0_121 br_0_121 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c121
*+ bl_0_121 br_0_121 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c121
*+ bl_0_121 br_0_121 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c121
*+ bl_0_121 br_0_121 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c121
*+ bl_0_121 br_0_121 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c121
*+ bl_0_121 br_0_121 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c121
*+ bl_0_121 br_0_121 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c121
*+ bl_0_121 br_0_121 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c121
*+ bl_0_121 br_0_121 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c121
*+ bl_0_121 br_0_121 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c121
*+ bl_0_121 br_0_121 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c121
*+ bl_0_121 br_0_121 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c121
*+ bl_0_121 br_0_121 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c121
*+ bl_0_121 br_0_121 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c121
*+ bl_0_121 br_0_121 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c121
*+ bl_0_121 br_0_121 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c121
*+ bl_0_121 br_0_121 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c121
*+ bl_0_121 br_0_121 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c121
*+ bl_0_121 br_0_121 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c121
*+ bl_0_121 br_0_121 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c121
*+ bl_0_121 br_0_121 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c121
*+ bl_0_121 br_0_121 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c121
*+ bl_0_121 br_0_121 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c121
*+ bl_0_121 br_0_121 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c121
*+ bl_0_121 br_0_121 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c121
*+ bl_0_121 br_0_121 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c121
*+ bl_0_121 br_0_121 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c121
*+ bl_0_121 br_0_121 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c121
*+ bl_0_121 br_0_121 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c121
*+ bl_0_121 br_0_121 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c121
*+ bl_0_121 br_0_121 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c121
*+ bl_0_121 br_0_121 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c121
*+ bl_0_121 br_0_121 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c121
*+ bl_0_121 br_0_121 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c121
*+ bl_0_121 br_0_121 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c121
*+ bl_0_121 br_0_121 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c121
*+ bl_0_121 br_0_121 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c121
*+ bl_0_121 br_0_121 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c121
*+ bl_0_121 br_0_121 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c121
*+ bl_0_121 br_0_121 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c121
*+ bl_0_121 br_0_121 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c121
*+ bl_0_121 br_0_121 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c121
*+ bl_0_121 br_0_121 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c121
*+ bl_0_121 br_0_121 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c121
*+ bl_0_121 br_0_121 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c121
*+ bl_0_121 br_0_121 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c121
*+ bl_0_121 br_0_121 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c121
*+ bl_0_121 br_0_121 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c121
*+ bl_0_121 br_0_121 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c121
*+ bl_0_121 br_0_121 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c121
*+ bl_0_121 br_0_121 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c121
*+ bl_0_121 br_0_121 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c121
*+ bl_0_121 br_0_121 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c121
*+ bl_0_121 br_0_121 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c121
*+ bl_0_121 br_0_121 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c121
*+ bl_0_121 br_0_121 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c121
*+ bl_0_121 br_0_121 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c121
*+ bl_0_121 br_0_121 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c121
*+ bl_0_121 br_0_121 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c121
*+ bl_0_121 br_0_121 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c121
*+ bl_0_121 br_0_121 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c121
*+ bl_0_121 br_0_121 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c121
*+ bl_0_121 br_0_121 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c121
*+ bl_0_121 br_0_121 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c121
*+ bl_0_121 br_0_121 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c121
*+ bl_0_121 br_0_121 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c121
*+ bl_0_121 br_0_121 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c121
*+ bl_0_121 br_0_121 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c121
*+ bl_0_121 br_0_121 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c121
*+ bl_0_121 br_0_121 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c121
*+ bl_0_121 br_0_121 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c121
*+ bl_0_121 br_0_121 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c121
*+ bl_0_121 br_0_121 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c121
*+ bl_0_121 br_0_121 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c121
*+ bl_0_121 br_0_121 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c121
*+ bl_0_121 br_0_121 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c121
*+ bl_0_121 br_0_121 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c121
*+ bl_0_121 br_0_121 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c121
*+ bl_0_121 br_0_121 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c121
*+ bl_0_121 br_0_121 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c121
*+ bl_0_121 br_0_121 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c121
*+ bl_0_121 br_0_121 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c121
*+ bl_0_121 br_0_121 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c121
*+ bl_0_121 br_0_121 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c121
*+ bl_0_121 br_0_121 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c121
*+ bl_0_121 br_0_121 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c121
*+ bl_0_121 br_0_121 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c121
*+ bl_0_121 br_0_121 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c121
*+ bl_0_121 br_0_121 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c121
*+ bl_0_121 br_0_121 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c121
*+ bl_0_121 br_0_121 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c121
*+ bl_0_121 br_0_121 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c121
*+ bl_0_121 br_0_121 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c121
*+ bl_0_121 br_0_121 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c121
*+ bl_0_121 br_0_121 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c121
*+ bl_0_121 br_0_121 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c121
*+ bl_0_121 br_0_121 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c121
*+ bl_0_121 br_0_121 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c121
*+ bl_0_121 br_0_121 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c121
*+ bl_0_121 br_0_121 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c121
*+ bl_0_121 br_0_121 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c121
*+ bl_0_121 br_0_121 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c121
*+ bl_0_121 br_0_121 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c121
*+ bl_0_121 br_0_121 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c121
*+ bl_0_121 br_0_121 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c121
*+ bl_0_121 br_0_121 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c121
*+ bl_0_121 br_0_121 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c121
*+ bl_0_121 br_0_121 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c121
*+ bl_0_121 br_0_121 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c121
*+ bl_0_121 br_0_121 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c121
*+ bl_0_121 br_0_121 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c121
*+ bl_0_121 br_0_121 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c121
*+ bl_0_121 br_0_121 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c121
*+ bl_0_121 br_0_121 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c121
*+ bl_0_121 br_0_121 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c121
*+ bl_0_121 br_0_121 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c121
*+ bl_0_121 br_0_121 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c121
*+ bl_0_121 br_0_121 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c121
*+ bl_0_121 br_0_121 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c121
*+ bl_0_121 br_0_121 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c121
*+ bl_0_121 br_0_121 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c121
*+ bl_0_121 br_0_121 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c121
*+ bl_0_121 br_0_121 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c121
*+ bl_0_121 br_0_121 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c121
*+ bl_0_121 br_0_121 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c121
*+ bl_0_121 br_0_121 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c121
+ bl_0_121 br_0_121 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c122
+ bl_0_122 br_0_122 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c122
*+ bl_0_122 br_0_122 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c122
*+ bl_0_122 br_0_122 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c122
*+ bl_0_122 br_0_122 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c122
*+ bl_0_122 br_0_122 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c122
*+ bl_0_122 br_0_122 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c122
*+ bl_0_122 br_0_122 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c122
*+ bl_0_122 br_0_122 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c122
*+ bl_0_122 br_0_122 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c122
*+ bl_0_122 br_0_122 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c122
*+ bl_0_122 br_0_122 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c122
*+ bl_0_122 br_0_122 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c122
*+ bl_0_122 br_0_122 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c122
*+ bl_0_122 br_0_122 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c122
*+ bl_0_122 br_0_122 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c122
*+ bl_0_122 br_0_122 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c122
*+ bl_0_122 br_0_122 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c122
*+ bl_0_122 br_0_122 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c122
*+ bl_0_122 br_0_122 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c122
*+ bl_0_122 br_0_122 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c122
*+ bl_0_122 br_0_122 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c122
*+ bl_0_122 br_0_122 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c122
*+ bl_0_122 br_0_122 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c122
*+ bl_0_122 br_0_122 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c122
*+ bl_0_122 br_0_122 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c122
*+ bl_0_122 br_0_122 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c122
*+ bl_0_122 br_0_122 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c122
*+ bl_0_122 br_0_122 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c122
*+ bl_0_122 br_0_122 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c122
*+ bl_0_122 br_0_122 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c122
*+ bl_0_122 br_0_122 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c122
*+ bl_0_122 br_0_122 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c122
*+ bl_0_122 br_0_122 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c122
*+ bl_0_122 br_0_122 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c122
*+ bl_0_122 br_0_122 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c122
*+ bl_0_122 br_0_122 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c122
*+ bl_0_122 br_0_122 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c122
*+ bl_0_122 br_0_122 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c122
*+ bl_0_122 br_0_122 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c122
*+ bl_0_122 br_0_122 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c122
*+ bl_0_122 br_0_122 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c122
*+ bl_0_122 br_0_122 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c122
*+ bl_0_122 br_0_122 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c122
*+ bl_0_122 br_0_122 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c122
*+ bl_0_122 br_0_122 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c122
*+ bl_0_122 br_0_122 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c122
*+ bl_0_122 br_0_122 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c122
*+ bl_0_122 br_0_122 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c122
*+ bl_0_122 br_0_122 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c122
*+ bl_0_122 br_0_122 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c122
*+ bl_0_122 br_0_122 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c122
*+ bl_0_122 br_0_122 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c122
*+ bl_0_122 br_0_122 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c122
*+ bl_0_122 br_0_122 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c122
*+ bl_0_122 br_0_122 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c122
*+ bl_0_122 br_0_122 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c122
*+ bl_0_122 br_0_122 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c122
*+ bl_0_122 br_0_122 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c122
*+ bl_0_122 br_0_122 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c122
*+ bl_0_122 br_0_122 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c122
*+ bl_0_122 br_0_122 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c122
*+ bl_0_122 br_0_122 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c122
*+ bl_0_122 br_0_122 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c122
*+ bl_0_122 br_0_122 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c122
*+ bl_0_122 br_0_122 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c122
*+ bl_0_122 br_0_122 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c122
*+ bl_0_122 br_0_122 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c122
*+ bl_0_122 br_0_122 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c122
*+ bl_0_122 br_0_122 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c122
*+ bl_0_122 br_0_122 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c122
*+ bl_0_122 br_0_122 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c122
*+ bl_0_122 br_0_122 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c122
*+ bl_0_122 br_0_122 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c122
*+ bl_0_122 br_0_122 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c122
*+ bl_0_122 br_0_122 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c122
*+ bl_0_122 br_0_122 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c122
*+ bl_0_122 br_0_122 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c122
*+ bl_0_122 br_0_122 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c122
*+ bl_0_122 br_0_122 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c122
*+ bl_0_122 br_0_122 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c122
*+ bl_0_122 br_0_122 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c122
*+ bl_0_122 br_0_122 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c122
*+ bl_0_122 br_0_122 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c122
*+ bl_0_122 br_0_122 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c122
*+ bl_0_122 br_0_122 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c122
*+ bl_0_122 br_0_122 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c122
*+ bl_0_122 br_0_122 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c122
*+ bl_0_122 br_0_122 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c122
*+ bl_0_122 br_0_122 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c122
*+ bl_0_122 br_0_122 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c122
*+ bl_0_122 br_0_122 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c122
*+ bl_0_122 br_0_122 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c122
*+ bl_0_122 br_0_122 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c122
*+ bl_0_122 br_0_122 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c122
*+ bl_0_122 br_0_122 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c122
*+ bl_0_122 br_0_122 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c122
*+ bl_0_122 br_0_122 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c122
*+ bl_0_122 br_0_122 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c122
*+ bl_0_122 br_0_122 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c122
*+ bl_0_122 br_0_122 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c122
*+ bl_0_122 br_0_122 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c122
*+ bl_0_122 br_0_122 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c122
*+ bl_0_122 br_0_122 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c122
*+ bl_0_122 br_0_122 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c122
*+ bl_0_122 br_0_122 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c122
*+ bl_0_122 br_0_122 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c122
*+ bl_0_122 br_0_122 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c122
*+ bl_0_122 br_0_122 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c122
*+ bl_0_122 br_0_122 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c122
*+ bl_0_122 br_0_122 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c122
*+ bl_0_122 br_0_122 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c122
*+ bl_0_122 br_0_122 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c122
*+ bl_0_122 br_0_122 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c122
*+ bl_0_122 br_0_122 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c122
*+ bl_0_122 br_0_122 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c122
*+ bl_0_122 br_0_122 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c122
*+ bl_0_122 br_0_122 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c122
*+ bl_0_122 br_0_122 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c122
*+ bl_0_122 br_0_122 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c122
*+ bl_0_122 br_0_122 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c122
*+ bl_0_122 br_0_122 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c122
*+ bl_0_122 br_0_122 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c122
*+ bl_0_122 br_0_122 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c122
*+ bl_0_122 br_0_122 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c122
*+ bl_0_122 br_0_122 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c122
*+ bl_0_122 br_0_122 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c122
*+ bl_0_122 br_0_122 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c122
+ bl_0_122 br_0_122 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c123
+ bl_0_123 br_0_123 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c123
*+ bl_0_123 br_0_123 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c123
*+ bl_0_123 br_0_123 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c123
*+ bl_0_123 br_0_123 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c123
*+ bl_0_123 br_0_123 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c123
*+ bl_0_123 br_0_123 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c123
*+ bl_0_123 br_0_123 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c123
*+ bl_0_123 br_0_123 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c123
*+ bl_0_123 br_0_123 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c123
*+ bl_0_123 br_0_123 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c123
*+ bl_0_123 br_0_123 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c123
*+ bl_0_123 br_0_123 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c123
*+ bl_0_123 br_0_123 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c123
*+ bl_0_123 br_0_123 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c123
*+ bl_0_123 br_0_123 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c123
*+ bl_0_123 br_0_123 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c123
*+ bl_0_123 br_0_123 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c123
*+ bl_0_123 br_0_123 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c123
*+ bl_0_123 br_0_123 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c123
*+ bl_0_123 br_0_123 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c123
*+ bl_0_123 br_0_123 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c123
*+ bl_0_123 br_0_123 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c123
*+ bl_0_123 br_0_123 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c123
*+ bl_0_123 br_0_123 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c123
*+ bl_0_123 br_0_123 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c123
*+ bl_0_123 br_0_123 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c123
*+ bl_0_123 br_0_123 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c123
*+ bl_0_123 br_0_123 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c123
*+ bl_0_123 br_0_123 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c123
*+ bl_0_123 br_0_123 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c123
*+ bl_0_123 br_0_123 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c123
*+ bl_0_123 br_0_123 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c123
*+ bl_0_123 br_0_123 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c123
*+ bl_0_123 br_0_123 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c123
*+ bl_0_123 br_0_123 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c123
*+ bl_0_123 br_0_123 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c123
*+ bl_0_123 br_0_123 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c123
*+ bl_0_123 br_0_123 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c123
*+ bl_0_123 br_0_123 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c123
*+ bl_0_123 br_0_123 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c123
*+ bl_0_123 br_0_123 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c123
*+ bl_0_123 br_0_123 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c123
*+ bl_0_123 br_0_123 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c123
*+ bl_0_123 br_0_123 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c123
*+ bl_0_123 br_0_123 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c123
*+ bl_0_123 br_0_123 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c123
*+ bl_0_123 br_0_123 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c123
*+ bl_0_123 br_0_123 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c123
*+ bl_0_123 br_0_123 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c123
*+ bl_0_123 br_0_123 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c123
*+ bl_0_123 br_0_123 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c123
*+ bl_0_123 br_0_123 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c123
*+ bl_0_123 br_0_123 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c123
*+ bl_0_123 br_0_123 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c123
*+ bl_0_123 br_0_123 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c123
*+ bl_0_123 br_0_123 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c123
*+ bl_0_123 br_0_123 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c123
*+ bl_0_123 br_0_123 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c123
*+ bl_0_123 br_0_123 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c123
*+ bl_0_123 br_0_123 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c123
*+ bl_0_123 br_0_123 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c123
*+ bl_0_123 br_0_123 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c123
*+ bl_0_123 br_0_123 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c123
*+ bl_0_123 br_0_123 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c123
*+ bl_0_123 br_0_123 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c123
*+ bl_0_123 br_0_123 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c123
*+ bl_0_123 br_0_123 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c123
*+ bl_0_123 br_0_123 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c123
*+ bl_0_123 br_0_123 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c123
*+ bl_0_123 br_0_123 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c123
*+ bl_0_123 br_0_123 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c123
*+ bl_0_123 br_0_123 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c123
*+ bl_0_123 br_0_123 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c123
*+ bl_0_123 br_0_123 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c123
*+ bl_0_123 br_0_123 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c123
*+ bl_0_123 br_0_123 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c123
*+ bl_0_123 br_0_123 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c123
*+ bl_0_123 br_0_123 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c123
*+ bl_0_123 br_0_123 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c123
*+ bl_0_123 br_0_123 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c123
*+ bl_0_123 br_0_123 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c123
*+ bl_0_123 br_0_123 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c123
*+ bl_0_123 br_0_123 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c123
*+ bl_0_123 br_0_123 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c123
*+ bl_0_123 br_0_123 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c123
*+ bl_0_123 br_0_123 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c123
*+ bl_0_123 br_0_123 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c123
*+ bl_0_123 br_0_123 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c123
*+ bl_0_123 br_0_123 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c123
*+ bl_0_123 br_0_123 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c123
*+ bl_0_123 br_0_123 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c123
*+ bl_0_123 br_0_123 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c123
*+ bl_0_123 br_0_123 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c123
*+ bl_0_123 br_0_123 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c123
*+ bl_0_123 br_0_123 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c123
*+ bl_0_123 br_0_123 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c123
*+ bl_0_123 br_0_123 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c123
*+ bl_0_123 br_0_123 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c123
*+ bl_0_123 br_0_123 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c123
*+ bl_0_123 br_0_123 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c123
*+ bl_0_123 br_0_123 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c123
*+ bl_0_123 br_0_123 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c123
*+ bl_0_123 br_0_123 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c123
*+ bl_0_123 br_0_123 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c123
*+ bl_0_123 br_0_123 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c123
*+ bl_0_123 br_0_123 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c123
*+ bl_0_123 br_0_123 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c123
*+ bl_0_123 br_0_123 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c123
*+ bl_0_123 br_0_123 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c123
*+ bl_0_123 br_0_123 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c123
*+ bl_0_123 br_0_123 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c123
*+ bl_0_123 br_0_123 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c123
*+ bl_0_123 br_0_123 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c123
*+ bl_0_123 br_0_123 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c123
*+ bl_0_123 br_0_123 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c123
*+ bl_0_123 br_0_123 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c123
*+ bl_0_123 br_0_123 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c123
*+ bl_0_123 br_0_123 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c123
*+ bl_0_123 br_0_123 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c123
*+ bl_0_123 br_0_123 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c123
*+ bl_0_123 br_0_123 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c123
*+ bl_0_123 br_0_123 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c123
*+ bl_0_123 br_0_123 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c123
*+ bl_0_123 br_0_123 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c123
*+ bl_0_123 br_0_123 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c123
*+ bl_0_123 br_0_123 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c123
*+ bl_0_123 br_0_123 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c123
+ bl_0_123 br_0_123 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c124
+ bl_0_124 br_0_124 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c124
*+ bl_0_124 br_0_124 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c124
*+ bl_0_124 br_0_124 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c124
*+ bl_0_124 br_0_124 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c124
*+ bl_0_124 br_0_124 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c124
*+ bl_0_124 br_0_124 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c124
*+ bl_0_124 br_0_124 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c124
*+ bl_0_124 br_0_124 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c124
*+ bl_0_124 br_0_124 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c124
*+ bl_0_124 br_0_124 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c124
*+ bl_0_124 br_0_124 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c124
*+ bl_0_124 br_0_124 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c124
*+ bl_0_124 br_0_124 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c124
*+ bl_0_124 br_0_124 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c124
*+ bl_0_124 br_0_124 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c124
*+ bl_0_124 br_0_124 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c124
*+ bl_0_124 br_0_124 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c124
*+ bl_0_124 br_0_124 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c124
*+ bl_0_124 br_0_124 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c124
*+ bl_0_124 br_0_124 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c124
*+ bl_0_124 br_0_124 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c124
*+ bl_0_124 br_0_124 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c124
*+ bl_0_124 br_0_124 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c124
*+ bl_0_124 br_0_124 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c124
*+ bl_0_124 br_0_124 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c124
*+ bl_0_124 br_0_124 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c124
*+ bl_0_124 br_0_124 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c124
*+ bl_0_124 br_0_124 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c124
*+ bl_0_124 br_0_124 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c124
*+ bl_0_124 br_0_124 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c124
*+ bl_0_124 br_0_124 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c124
*+ bl_0_124 br_0_124 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c124
*+ bl_0_124 br_0_124 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c124
*+ bl_0_124 br_0_124 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c124
*+ bl_0_124 br_0_124 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c124
*+ bl_0_124 br_0_124 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c124
*+ bl_0_124 br_0_124 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c124
*+ bl_0_124 br_0_124 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c124
*+ bl_0_124 br_0_124 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c124
*+ bl_0_124 br_0_124 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c124
*+ bl_0_124 br_0_124 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c124
*+ bl_0_124 br_0_124 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c124
*+ bl_0_124 br_0_124 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c124
*+ bl_0_124 br_0_124 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c124
*+ bl_0_124 br_0_124 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c124
*+ bl_0_124 br_0_124 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c124
*+ bl_0_124 br_0_124 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c124
*+ bl_0_124 br_0_124 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c124
*+ bl_0_124 br_0_124 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c124
*+ bl_0_124 br_0_124 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c124
*+ bl_0_124 br_0_124 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c124
*+ bl_0_124 br_0_124 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c124
*+ bl_0_124 br_0_124 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c124
*+ bl_0_124 br_0_124 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c124
*+ bl_0_124 br_0_124 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c124
*+ bl_0_124 br_0_124 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c124
*+ bl_0_124 br_0_124 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c124
*+ bl_0_124 br_0_124 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c124
*+ bl_0_124 br_0_124 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c124
*+ bl_0_124 br_0_124 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c124
*+ bl_0_124 br_0_124 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c124
*+ bl_0_124 br_0_124 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c124
*+ bl_0_124 br_0_124 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c124
*+ bl_0_124 br_0_124 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c124
*+ bl_0_124 br_0_124 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c124
*+ bl_0_124 br_0_124 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c124
*+ bl_0_124 br_0_124 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c124
*+ bl_0_124 br_0_124 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c124
*+ bl_0_124 br_0_124 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c124
*+ bl_0_124 br_0_124 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c124
*+ bl_0_124 br_0_124 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c124
*+ bl_0_124 br_0_124 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c124
*+ bl_0_124 br_0_124 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c124
*+ bl_0_124 br_0_124 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c124
*+ bl_0_124 br_0_124 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c124
*+ bl_0_124 br_0_124 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c124
*+ bl_0_124 br_0_124 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c124
*+ bl_0_124 br_0_124 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c124
*+ bl_0_124 br_0_124 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c124
*+ bl_0_124 br_0_124 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c124
*+ bl_0_124 br_0_124 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c124
*+ bl_0_124 br_0_124 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c124
*+ bl_0_124 br_0_124 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c124
*+ bl_0_124 br_0_124 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c124
*+ bl_0_124 br_0_124 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c124
*+ bl_0_124 br_0_124 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c124
*+ bl_0_124 br_0_124 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c124
*+ bl_0_124 br_0_124 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c124
*+ bl_0_124 br_0_124 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c124
*+ bl_0_124 br_0_124 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c124
*+ bl_0_124 br_0_124 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c124
*+ bl_0_124 br_0_124 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c124
*+ bl_0_124 br_0_124 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c124
*+ bl_0_124 br_0_124 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c124
*+ bl_0_124 br_0_124 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c124
*+ bl_0_124 br_0_124 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c124
*+ bl_0_124 br_0_124 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c124
*+ bl_0_124 br_0_124 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c124
*+ bl_0_124 br_0_124 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c124
*+ bl_0_124 br_0_124 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c124
*+ bl_0_124 br_0_124 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c124
*+ bl_0_124 br_0_124 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c124
*+ bl_0_124 br_0_124 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c124
*+ bl_0_124 br_0_124 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c124
*+ bl_0_124 br_0_124 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c124
*+ bl_0_124 br_0_124 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c124
*+ bl_0_124 br_0_124 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c124
*+ bl_0_124 br_0_124 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c124
*+ bl_0_124 br_0_124 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c124
*+ bl_0_124 br_0_124 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c124
*+ bl_0_124 br_0_124 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c124
*+ bl_0_124 br_0_124 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c124
*+ bl_0_124 br_0_124 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c124
*+ bl_0_124 br_0_124 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c124
*+ bl_0_124 br_0_124 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c124
*+ bl_0_124 br_0_124 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c124
*+ bl_0_124 br_0_124 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c124
*+ bl_0_124 br_0_124 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c124
*+ bl_0_124 br_0_124 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c124
*+ bl_0_124 br_0_124 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c124
*+ bl_0_124 br_0_124 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c124
*+ bl_0_124 br_0_124 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c124
*+ bl_0_124 br_0_124 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c124
*+ bl_0_124 br_0_124 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c124
*+ bl_0_124 br_0_124 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c124
*+ bl_0_124 br_0_124 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c124
*+ bl_0_124 br_0_124 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c124
+ bl_0_124 br_0_124 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c125
+ bl_0_125 br_0_125 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c125
*+ bl_0_125 br_0_125 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c125
*+ bl_0_125 br_0_125 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c125
*+ bl_0_125 br_0_125 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c125
*+ bl_0_125 br_0_125 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c125
*+ bl_0_125 br_0_125 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c125
*+ bl_0_125 br_0_125 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c125
*+ bl_0_125 br_0_125 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c125
*+ bl_0_125 br_0_125 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c125
*+ bl_0_125 br_0_125 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c125
*+ bl_0_125 br_0_125 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c125
*+ bl_0_125 br_0_125 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c125
*+ bl_0_125 br_0_125 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c125
*+ bl_0_125 br_0_125 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c125
*+ bl_0_125 br_0_125 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c125
*+ bl_0_125 br_0_125 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c125
*+ bl_0_125 br_0_125 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c125
*+ bl_0_125 br_0_125 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c125
*+ bl_0_125 br_0_125 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c125
*+ bl_0_125 br_0_125 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c125
*+ bl_0_125 br_0_125 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c125
*+ bl_0_125 br_0_125 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c125
*+ bl_0_125 br_0_125 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c125
*+ bl_0_125 br_0_125 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c125
*+ bl_0_125 br_0_125 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c125
*+ bl_0_125 br_0_125 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c125
*+ bl_0_125 br_0_125 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c125
*+ bl_0_125 br_0_125 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c125
*+ bl_0_125 br_0_125 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c125
*+ bl_0_125 br_0_125 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c125
*+ bl_0_125 br_0_125 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c125
*+ bl_0_125 br_0_125 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c125
*+ bl_0_125 br_0_125 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c125
*+ bl_0_125 br_0_125 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c125
*+ bl_0_125 br_0_125 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c125
*+ bl_0_125 br_0_125 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c125
*+ bl_0_125 br_0_125 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c125
*+ bl_0_125 br_0_125 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c125
*+ bl_0_125 br_0_125 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c125
*+ bl_0_125 br_0_125 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c125
*+ bl_0_125 br_0_125 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c125
*+ bl_0_125 br_0_125 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c125
*+ bl_0_125 br_0_125 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c125
*+ bl_0_125 br_0_125 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c125
*+ bl_0_125 br_0_125 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c125
*+ bl_0_125 br_0_125 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c125
*+ bl_0_125 br_0_125 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c125
*+ bl_0_125 br_0_125 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c125
*+ bl_0_125 br_0_125 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c125
*+ bl_0_125 br_0_125 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c125
*+ bl_0_125 br_0_125 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c125
*+ bl_0_125 br_0_125 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c125
*+ bl_0_125 br_0_125 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c125
*+ bl_0_125 br_0_125 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c125
*+ bl_0_125 br_0_125 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c125
*+ bl_0_125 br_0_125 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c125
*+ bl_0_125 br_0_125 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c125
*+ bl_0_125 br_0_125 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c125
*+ bl_0_125 br_0_125 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c125
*+ bl_0_125 br_0_125 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c125
*+ bl_0_125 br_0_125 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c125
*+ bl_0_125 br_0_125 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c125
*+ bl_0_125 br_0_125 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c125
*+ bl_0_125 br_0_125 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c125
*+ bl_0_125 br_0_125 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c125
*+ bl_0_125 br_0_125 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c125
*+ bl_0_125 br_0_125 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c125
*+ bl_0_125 br_0_125 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c125
*+ bl_0_125 br_0_125 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c125
*+ bl_0_125 br_0_125 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c125
*+ bl_0_125 br_0_125 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c125
*+ bl_0_125 br_0_125 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c125
*+ bl_0_125 br_0_125 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c125
*+ bl_0_125 br_0_125 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c125
*+ bl_0_125 br_0_125 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c125
*+ bl_0_125 br_0_125 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c125
*+ bl_0_125 br_0_125 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c125
*+ bl_0_125 br_0_125 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c125
*+ bl_0_125 br_0_125 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c125
*+ bl_0_125 br_0_125 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c125
*+ bl_0_125 br_0_125 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c125
*+ bl_0_125 br_0_125 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c125
*+ bl_0_125 br_0_125 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c125
*+ bl_0_125 br_0_125 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c125
*+ bl_0_125 br_0_125 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c125
*+ bl_0_125 br_0_125 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c125
*+ bl_0_125 br_0_125 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c125
*+ bl_0_125 br_0_125 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c125
*+ bl_0_125 br_0_125 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c125
*+ bl_0_125 br_0_125 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c125
*+ bl_0_125 br_0_125 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c125
*+ bl_0_125 br_0_125 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c125
*+ bl_0_125 br_0_125 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c125
*+ bl_0_125 br_0_125 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c125
*+ bl_0_125 br_0_125 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c125
*+ bl_0_125 br_0_125 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c125
*+ bl_0_125 br_0_125 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c125
*+ bl_0_125 br_0_125 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c125
*+ bl_0_125 br_0_125 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c125
*+ bl_0_125 br_0_125 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c125
*+ bl_0_125 br_0_125 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c125
*+ bl_0_125 br_0_125 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c125
*+ bl_0_125 br_0_125 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c125
*+ bl_0_125 br_0_125 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c125
*+ bl_0_125 br_0_125 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c125
*+ bl_0_125 br_0_125 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c125
*+ bl_0_125 br_0_125 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c125
*+ bl_0_125 br_0_125 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c125
*+ bl_0_125 br_0_125 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c125
*+ bl_0_125 br_0_125 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c125
*+ bl_0_125 br_0_125 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c125
*+ bl_0_125 br_0_125 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c125
*+ bl_0_125 br_0_125 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c125
*+ bl_0_125 br_0_125 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c125
*+ bl_0_125 br_0_125 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c125
*+ bl_0_125 br_0_125 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c125
*+ bl_0_125 br_0_125 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c125
*+ bl_0_125 br_0_125 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c125
*+ bl_0_125 br_0_125 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c125
*+ bl_0_125 br_0_125 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c125
*+ bl_0_125 br_0_125 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c125
*+ bl_0_125 br_0_125 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c125
*+ bl_0_125 br_0_125 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c125
*+ bl_0_125 br_0_125 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c125
*+ bl_0_125 br_0_125 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c125
*+ bl_0_125 br_0_125 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c125
*+ bl_0_125 br_0_125 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c125
+ bl_0_125 br_0_125 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c126
+ bl_0_126 br_0_126 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c126
*+ bl_0_126 br_0_126 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c126
*+ bl_0_126 br_0_126 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c126
*+ bl_0_126 br_0_126 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c126
*+ bl_0_126 br_0_126 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c126
*+ bl_0_126 br_0_126 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c126
*+ bl_0_126 br_0_126 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c126
*+ bl_0_126 br_0_126 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c126
*+ bl_0_126 br_0_126 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c126
*+ bl_0_126 br_0_126 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c126
*+ bl_0_126 br_0_126 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c126
*+ bl_0_126 br_0_126 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c126
*+ bl_0_126 br_0_126 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c126
*+ bl_0_126 br_0_126 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c126
*+ bl_0_126 br_0_126 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c126
*+ bl_0_126 br_0_126 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c126
*+ bl_0_126 br_0_126 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c126
*+ bl_0_126 br_0_126 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c126
*+ bl_0_126 br_0_126 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c126
*+ bl_0_126 br_0_126 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c126
*+ bl_0_126 br_0_126 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c126
*+ bl_0_126 br_0_126 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c126
*+ bl_0_126 br_0_126 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c126
*+ bl_0_126 br_0_126 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c126
*+ bl_0_126 br_0_126 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c126
*+ bl_0_126 br_0_126 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c126
*+ bl_0_126 br_0_126 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c126
*+ bl_0_126 br_0_126 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c126
*+ bl_0_126 br_0_126 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c126
*+ bl_0_126 br_0_126 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c126
*+ bl_0_126 br_0_126 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c126
*+ bl_0_126 br_0_126 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c126
*+ bl_0_126 br_0_126 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c126
*+ bl_0_126 br_0_126 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c126
*+ bl_0_126 br_0_126 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c126
*+ bl_0_126 br_0_126 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c126
*+ bl_0_126 br_0_126 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c126
*+ bl_0_126 br_0_126 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c126
*+ bl_0_126 br_0_126 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c126
*+ bl_0_126 br_0_126 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c126
*+ bl_0_126 br_0_126 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c126
*+ bl_0_126 br_0_126 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c126
*+ bl_0_126 br_0_126 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c126
*+ bl_0_126 br_0_126 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c126
*+ bl_0_126 br_0_126 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c126
*+ bl_0_126 br_0_126 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c126
*+ bl_0_126 br_0_126 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c126
*+ bl_0_126 br_0_126 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c126
*+ bl_0_126 br_0_126 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c126
*+ bl_0_126 br_0_126 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c126
*+ bl_0_126 br_0_126 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c126
*+ bl_0_126 br_0_126 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c126
*+ bl_0_126 br_0_126 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c126
*+ bl_0_126 br_0_126 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c126
*+ bl_0_126 br_0_126 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c126
*+ bl_0_126 br_0_126 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c126
*+ bl_0_126 br_0_126 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c126
*+ bl_0_126 br_0_126 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c126
*+ bl_0_126 br_0_126 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c126
*+ bl_0_126 br_0_126 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c126
*+ bl_0_126 br_0_126 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c126
*+ bl_0_126 br_0_126 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c126
*+ bl_0_126 br_0_126 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c126
*+ bl_0_126 br_0_126 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c126
*+ bl_0_126 br_0_126 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c126
*+ bl_0_126 br_0_126 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c126
*+ bl_0_126 br_0_126 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c126
*+ bl_0_126 br_0_126 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c126
*+ bl_0_126 br_0_126 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c126
*+ bl_0_126 br_0_126 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c126
*+ bl_0_126 br_0_126 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c126
*+ bl_0_126 br_0_126 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c126
*+ bl_0_126 br_0_126 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c126
*+ bl_0_126 br_0_126 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c126
*+ bl_0_126 br_0_126 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c126
*+ bl_0_126 br_0_126 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c126
*+ bl_0_126 br_0_126 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c126
*+ bl_0_126 br_0_126 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c126
*+ bl_0_126 br_0_126 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c126
*+ bl_0_126 br_0_126 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c126
*+ bl_0_126 br_0_126 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c126
*+ bl_0_126 br_0_126 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c126
*+ bl_0_126 br_0_126 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c126
*+ bl_0_126 br_0_126 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c126
*+ bl_0_126 br_0_126 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c126
*+ bl_0_126 br_0_126 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c126
*+ bl_0_126 br_0_126 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c126
*+ bl_0_126 br_0_126 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c126
*+ bl_0_126 br_0_126 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c126
*+ bl_0_126 br_0_126 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c126
*+ bl_0_126 br_0_126 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c126
*+ bl_0_126 br_0_126 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c126
*+ bl_0_126 br_0_126 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c126
*+ bl_0_126 br_0_126 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c126
*+ bl_0_126 br_0_126 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c126
*+ bl_0_126 br_0_126 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c126
*+ bl_0_126 br_0_126 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c126
*+ bl_0_126 br_0_126 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c126
*+ bl_0_126 br_0_126 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c126
*+ bl_0_126 br_0_126 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c126
*+ bl_0_126 br_0_126 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c126
*+ bl_0_126 br_0_126 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c126
*+ bl_0_126 br_0_126 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c126
*+ bl_0_126 br_0_126 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c126
*+ bl_0_126 br_0_126 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c126
*+ bl_0_126 br_0_126 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c126
*+ bl_0_126 br_0_126 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c126
*+ bl_0_126 br_0_126 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c126
*+ bl_0_126 br_0_126 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c126
*+ bl_0_126 br_0_126 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c126
*+ bl_0_126 br_0_126 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c126
*+ bl_0_126 br_0_126 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c126
*+ bl_0_126 br_0_126 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c126
*+ bl_0_126 br_0_126 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c126
*+ bl_0_126 br_0_126 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c126
*+ bl_0_126 br_0_126 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c126
*+ bl_0_126 br_0_126 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c126
*+ bl_0_126 br_0_126 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c126
*+ bl_0_126 br_0_126 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c126
*+ bl_0_126 br_0_126 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c126
*+ bl_0_126 br_0_126 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c126
*+ bl_0_126 br_0_126 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c126
*+ bl_0_126 br_0_126 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c126
*+ bl_0_126 br_0_126 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c126
*+ bl_0_126 br_0_126 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c126
*+ bl_0_126 br_0_126 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c126
*+ bl_0_126 br_0_126 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c126
+ bl_0_126 br_0_126 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c127
+ bl_0_127 br_0_127 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c127
*+ bl_0_127 br_0_127 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c127
*+ bl_0_127 br_0_127 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c127
*+ bl_0_127 br_0_127 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c127
*+ bl_0_127 br_0_127 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c127
*+ bl_0_127 br_0_127 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c127
*+ bl_0_127 br_0_127 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c127
*+ bl_0_127 br_0_127 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c127
*+ bl_0_127 br_0_127 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c127
*+ bl_0_127 br_0_127 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c127
*+ bl_0_127 br_0_127 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c127
*+ bl_0_127 br_0_127 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c127
*+ bl_0_127 br_0_127 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c127
*+ bl_0_127 br_0_127 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c127
*+ bl_0_127 br_0_127 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c127
*+ bl_0_127 br_0_127 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c127
*+ bl_0_127 br_0_127 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c127
*+ bl_0_127 br_0_127 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c127
*+ bl_0_127 br_0_127 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c127
*+ bl_0_127 br_0_127 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c127
*+ bl_0_127 br_0_127 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c127
*+ bl_0_127 br_0_127 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c127
*+ bl_0_127 br_0_127 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c127
*+ bl_0_127 br_0_127 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c127
*+ bl_0_127 br_0_127 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c127
*+ bl_0_127 br_0_127 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c127
*+ bl_0_127 br_0_127 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c127
*+ bl_0_127 br_0_127 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c127
*+ bl_0_127 br_0_127 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c127
*+ bl_0_127 br_0_127 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c127
*+ bl_0_127 br_0_127 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c127
*+ bl_0_127 br_0_127 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c127
*+ bl_0_127 br_0_127 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c127
*+ bl_0_127 br_0_127 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c127
*+ bl_0_127 br_0_127 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c127
*+ bl_0_127 br_0_127 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c127
*+ bl_0_127 br_0_127 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c127
*+ bl_0_127 br_0_127 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c127
*+ bl_0_127 br_0_127 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c127
*+ bl_0_127 br_0_127 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c127
*+ bl_0_127 br_0_127 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c127
*+ bl_0_127 br_0_127 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c127
*+ bl_0_127 br_0_127 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c127
*+ bl_0_127 br_0_127 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c127
*+ bl_0_127 br_0_127 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c127
*+ bl_0_127 br_0_127 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c127
*+ bl_0_127 br_0_127 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c127
*+ bl_0_127 br_0_127 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c127
*+ bl_0_127 br_0_127 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c127
*+ bl_0_127 br_0_127 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c127
*+ bl_0_127 br_0_127 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c127
*+ bl_0_127 br_0_127 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c127
*+ bl_0_127 br_0_127 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c127
*+ bl_0_127 br_0_127 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c127
*+ bl_0_127 br_0_127 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c127
*+ bl_0_127 br_0_127 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c127
*+ bl_0_127 br_0_127 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c127
*+ bl_0_127 br_0_127 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c127
*+ bl_0_127 br_0_127 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c127
*+ bl_0_127 br_0_127 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c127
*+ bl_0_127 br_0_127 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c127
*+ bl_0_127 br_0_127 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c127
*+ bl_0_127 br_0_127 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c127
*+ bl_0_127 br_0_127 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c127
*+ bl_0_127 br_0_127 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c127
*+ bl_0_127 br_0_127 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c127
*+ bl_0_127 br_0_127 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c127
*+ bl_0_127 br_0_127 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c127
*+ bl_0_127 br_0_127 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c127
*+ bl_0_127 br_0_127 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c127
*+ bl_0_127 br_0_127 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c127
*+ bl_0_127 br_0_127 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c127
*+ bl_0_127 br_0_127 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c127
*+ bl_0_127 br_0_127 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c127
*+ bl_0_127 br_0_127 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c127
*+ bl_0_127 br_0_127 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c127
*+ bl_0_127 br_0_127 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c127
*+ bl_0_127 br_0_127 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c127
*+ bl_0_127 br_0_127 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c127
*+ bl_0_127 br_0_127 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c127
*+ bl_0_127 br_0_127 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c127
*+ bl_0_127 br_0_127 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c127
*+ bl_0_127 br_0_127 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c127
*+ bl_0_127 br_0_127 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c127
*+ bl_0_127 br_0_127 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c127
*+ bl_0_127 br_0_127 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c127
*+ bl_0_127 br_0_127 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c127
*+ bl_0_127 br_0_127 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c127
*+ bl_0_127 br_0_127 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c127
*+ bl_0_127 br_0_127 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c127
*+ bl_0_127 br_0_127 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c127
*+ bl_0_127 br_0_127 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c127
*+ bl_0_127 br_0_127 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c127
*+ bl_0_127 br_0_127 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c127
*+ bl_0_127 br_0_127 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c127
*+ bl_0_127 br_0_127 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c127
*+ bl_0_127 br_0_127 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c127
*+ bl_0_127 br_0_127 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c127
*+ bl_0_127 br_0_127 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c127
*+ bl_0_127 br_0_127 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c127
*+ bl_0_127 br_0_127 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c127
*+ bl_0_127 br_0_127 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c127
*+ bl_0_127 br_0_127 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c127
*+ bl_0_127 br_0_127 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c127
*+ bl_0_127 br_0_127 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c127
*+ bl_0_127 br_0_127 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c127
*+ bl_0_127 br_0_127 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c127
*+ bl_0_127 br_0_127 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c127
*+ bl_0_127 br_0_127 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c127
*+ bl_0_127 br_0_127 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c127
*+ bl_0_127 br_0_127 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c127
*+ bl_0_127 br_0_127 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c127
*+ bl_0_127 br_0_127 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c127
*+ bl_0_127 br_0_127 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c127
*+ bl_0_127 br_0_127 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c127
*+ bl_0_127 br_0_127 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c127
*+ bl_0_127 br_0_127 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c127
*+ bl_0_127 br_0_127 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c127
*+ bl_0_127 br_0_127 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c127
*+ bl_0_127 br_0_127 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c127
*+ bl_0_127 br_0_127 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c127
*+ bl_0_127 br_0_127 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c127
*+ bl_0_127 br_0_127 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c127
*+ bl_0_127 br_0_127 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c127
*+ bl_0_127 br_0_127 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c127
*+ bl_0_127 br_0_127 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c127
*+ bl_0_127 br_0_127 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c127
+ bl_0_127 br_0_127 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c128
+ bl_0_128 br_0_128 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c128
*+ bl_0_128 br_0_128 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c128
*+ bl_0_128 br_0_128 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c128
*+ bl_0_128 br_0_128 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c128
*+ bl_0_128 br_0_128 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c128
*+ bl_0_128 br_0_128 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c128
*+ bl_0_128 br_0_128 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c128
*+ bl_0_128 br_0_128 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c128
*+ bl_0_128 br_0_128 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c128
*+ bl_0_128 br_0_128 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c128
*+ bl_0_128 br_0_128 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c128
*+ bl_0_128 br_0_128 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c128
*+ bl_0_128 br_0_128 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c128
*+ bl_0_128 br_0_128 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c128
*+ bl_0_128 br_0_128 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c128
*+ bl_0_128 br_0_128 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c128
*+ bl_0_128 br_0_128 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c128
*+ bl_0_128 br_0_128 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c128
*+ bl_0_128 br_0_128 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c128
*+ bl_0_128 br_0_128 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c128
*+ bl_0_128 br_0_128 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c128
*+ bl_0_128 br_0_128 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c128
*+ bl_0_128 br_0_128 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c128
*+ bl_0_128 br_0_128 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c128
*+ bl_0_128 br_0_128 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c128
*+ bl_0_128 br_0_128 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c128
*+ bl_0_128 br_0_128 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c128
*+ bl_0_128 br_0_128 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c128
*+ bl_0_128 br_0_128 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c128
*+ bl_0_128 br_0_128 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c128
*+ bl_0_128 br_0_128 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c128
*+ bl_0_128 br_0_128 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c128
*+ bl_0_128 br_0_128 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c128
*+ bl_0_128 br_0_128 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c128
*+ bl_0_128 br_0_128 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c128
*+ bl_0_128 br_0_128 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c128
*+ bl_0_128 br_0_128 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c128
*+ bl_0_128 br_0_128 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c128
*+ bl_0_128 br_0_128 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c128
*+ bl_0_128 br_0_128 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c128
*+ bl_0_128 br_0_128 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c128
*+ bl_0_128 br_0_128 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c128
*+ bl_0_128 br_0_128 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c128
*+ bl_0_128 br_0_128 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c128
*+ bl_0_128 br_0_128 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c128
*+ bl_0_128 br_0_128 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c128
*+ bl_0_128 br_0_128 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c128
*+ bl_0_128 br_0_128 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c128
*+ bl_0_128 br_0_128 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c128
*+ bl_0_128 br_0_128 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c128
*+ bl_0_128 br_0_128 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c128
*+ bl_0_128 br_0_128 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c128
*+ bl_0_128 br_0_128 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c128
*+ bl_0_128 br_0_128 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c128
*+ bl_0_128 br_0_128 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c128
*+ bl_0_128 br_0_128 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c128
*+ bl_0_128 br_0_128 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c128
*+ bl_0_128 br_0_128 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c128
*+ bl_0_128 br_0_128 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c128
*+ bl_0_128 br_0_128 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c128
*+ bl_0_128 br_0_128 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c128
*+ bl_0_128 br_0_128 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c128
*+ bl_0_128 br_0_128 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c128
*+ bl_0_128 br_0_128 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c128
*+ bl_0_128 br_0_128 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c128
*+ bl_0_128 br_0_128 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c128
*+ bl_0_128 br_0_128 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c128
*+ bl_0_128 br_0_128 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c128
*+ bl_0_128 br_0_128 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c128
*+ bl_0_128 br_0_128 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c128
*+ bl_0_128 br_0_128 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c128
*+ bl_0_128 br_0_128 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c128
*+ bl_0_128 br_0_128 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c128
*+ bl_0_128 br_0_128 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c128
*+ bl_0_128 br_0_128 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c128
*+ bl_0_128 br_0_128 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c128
*+ bl_0_128 br_0_128 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c128
*+ bl_0_128 br_0_128 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c128
*+ bl_0_128 br_0_128 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c128
*+ bl_0_128 br_0_128 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c128
*+ bl_0_128 br_0_128 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c128
*+ bl_0_128 br_0_128 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c128
*+ bl_0_128 br_0_128 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c128
*+ bl_0_128 br_0_128 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c128
*+ bl_0_128 br_0_128 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c128
*+ bl_0_128 br_0_128 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c128
*+ bl_0_128 br_0_128 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c128
*+ bl_0_128 br_0_128 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c128
*+ bl_0_128 br_0_128 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c128
*+ bl_0_128 br_0_128 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c128
*+ bl_0_128 br_0_128 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c128
*+ bl_0_128 br_0_128 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c128
*+ bl_0_128 br_0_128 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c128
*+ bl_0_128 br_0_128 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c128
*+ bl_0_128 br_0_128 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c128
*+ bl_0_128 br_0_128 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c128
*+ bl_0_128 br_0_128 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c128
*+ bl_0_128 br_0_128 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c128
*+ bl_0_128 br_0_128 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c128
*+ bl_0_128 br_0_128 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c128
*+ bl_0_128 br_0_128 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c128
*+ bl_0_128 br_0_128 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c128
*+ bl_0_128 br_0_128 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c128
*+ bl_0_128 br_0_128 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c128
*+ bl_0_128 br_0_128 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c128
*+ bl_0_128 br_0_128 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c128
*+ bl_0_128 br_0_128 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c128
*+ bl_0_128 br_0_128 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c128
*+ bl_0_128 br_0_128 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c128
*+ bl_0_128 br_0_128 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c128
*+ bl_0_128 br_0_128 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c128
*+ bl_0_128 br_0_128 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c128
*+ bl_0_128 br_0_128 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c128
*+ bl_0_128 br_0_128 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c128
*+ bl_0_128 br_0_128 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c128
*+ bl_0_128 br_0_128 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c128
*+ bl_0_128 br_0_128 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c128
*+ bl_0_128 br_0_128 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c128
*+ bl_0_128 br_0_128 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c128
*+ bl_0_128 br_0_128 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c128
*+ bl_0_128 br_0_128 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c128
*+ bl_0_128 br_0_128 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c128
*+ bl_0_128 br_0_128 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c128
*+ bl_0_128 br_0_128 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c128
*+ bl_0_128 br_0_128 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c128
*+ bl_0_128 br_0_128 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c128
*+ bl_0_128 br_0_128 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c128
+ bl_0_128 br_0_128 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c129
+ bl_0_129 br_0_129 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c129
*+ bl_0_129 br_0_129 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c129
*+ bl_0_129 br_0_129 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c129
*+ bl_0_129 br_0_129 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c129
*+ bl_0_129 br_0_129 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c129
*+ bl_0_129 br_0_129 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c129
*+ bl_0_129 br_0_129 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c129
*+ bl_0_129 br_0_129 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c129
*+ bl_0_129 br_0_129 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c129
*+ bl_0_129 br_0_129 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c129
*+ bl_0_129 br_0_129 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c129
*+ bl_0_129 br_0_129 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c129
*+ bl_0_129 br_0_129 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c129
*+ bl_0_129 br_0_129 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c129
*+ bl_0_129 br_0_129 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c129
*+ bl_0_129 br_0_129 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c129
*+ bl_0_129 br_0_129 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c129
*+ bl_0_129 br_0_129 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c129
*+ bl_0_129 br_0_129 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c129
*+ bl_0_129 br_0_129 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c129
*+ bl_0_129 br_0_129 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c129
*+ bl_0_129 br_0_129 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c129
*+ bl_0_129 br_0_129 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c129
*+ bl_0_129 br_0_129 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c129
*+ bl_0_129 br_0_129 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c129
*+ bl_0_129 br_0_129 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c129
*+ bl_0_129 br_0_129 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c129
*+ bl_0_129 br_0_129 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c129
*+ bl_0_129 br_0_129 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c129
*+ bl_0_129 br_0_129 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c129
*+ bl_0_129 br_0_129 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c129
*+ bl_0_129 br_0_129 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c129
*+ bl_0_129 br_0_129 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c129
*+ bl_0_129 br_0_129 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c129
*+ bl_0_129 br_0_129 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c129
*+ bl_0_129 br_0_129 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c129
*+ bl_0_129 br_0_129 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c129
*+ bl_0_129 br_0_129 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c129
*+ bl_0_129 br_0_129 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c129
*+ bl_0_129 br_0_129 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c129
*+ bl_0_129 br_0_129 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c129
*+ bl_0_129 br_0_129 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c129
*+ bl_0_129 br_0_129 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c129
*+ bl_0_129 br_0_129 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c129
*+ bl_0_129 br_0_129 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c129
*+ bl_0_129 br_0_129 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c129
*+ bl_0_129 br_0_129 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c129
*+ bl_0_129 br_0_129 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c129
*+ bl_0_129 br_0_129 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c129
*+ bl_0_129 br_0_129 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c129
*+ bl_0_129 br_0_129 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c129
*+ bl_0_129 br_0_129 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c129
*+ bl_0_129 br_0_129 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c129
*+ bl_0_129 br_0_129 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c129
*+ bl_0_129 br_0_129 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c129
*+ bl_0_129 br_0_129 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c129
*+ bl_0_129 br_0_129 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c129
*+ bl_0_129 br_0_129 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c129
*+ bl_0_129 br_0_129 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c129
*+ bl_0_129 br_0_129 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c129
*+ bl_0_129 br_0_129 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c129
*+ bl_0_129 br_0_129 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c129
*+ bl_0_129 br_0_129 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c129
*+ bl_0_129 br_0_129 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c129
*+ bl_0_129 br_0_129 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c129
*+ bl_0_129 br_0_129 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c129
*+ bl_0_129 br_0_129 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c129
*+ bl_0_129 br_0_129 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c129
*+ bl_0_129 br_0_129 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c129
*+ bl_0_129 br_0_129 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c129
*+ bl_0_129 br_0_129 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c129
*+ bl_0_129 br_0_129 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c129
*+ bl_0_129 br_0_129 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c129
*+ bl_0_129 br_0_129 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c129
*+ bl_0_129 br_0_129 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c129
*+ bl_0_129 br_0_129 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c129
*+ bl_0_129 br_0_129 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c129
*+ bl_0_129 br_0_129 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c129
*+ bl_0_129 br_0_129 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c129
*+ bl_0_129 br_0_129 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c129
*+ bl_0_129 br_0_129 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c129
*+ bl_0_129 br_0_129 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c129
*+ bl_0_129 br_0_129 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c129
*+ bl_0_129 br_0_129 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c129
*+ bl_0_129 br_0_129 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c129
*+ bl_0_129 br_0_129 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c129
*+ bl_0_129 br_0_129 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c129
*+ bl_0_129 br_0_129 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c129
*+ bl_0_129 br_0_129 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c129
*+ bl_0_129 br_0_129 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c129
*+ bl_0_129 br_0_129 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c129
*+ bl_0_129 br_0_129 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c129
*+ bl_0_129 br_0_129 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c129
*+ bl_0_129 br_0_129 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c129
*+ bl_0_129 br_0_129 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c129
*+ bl_0_129 br_0_129 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c129
*+ bl_0_129 br_0_129 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c129
*+ bl_0_129 br_0_129 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c129
*+ bl_0_129 br_0_129 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c129
*+ bl_0_129 br_0_129 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c129
*+ bl_0_129 br_0_129 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c129
*+ bl_0_129 br_0_129 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c129
*+ bl_0_129 br_0_129 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c129
*+ bl_0_129 br_0_129 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c129
*+ bl_0_129 br_0_129 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c129
*+ bl_0_129 br_0_129 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c129
*+ bl_0_129 br_0_129 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c129
*+ bl_0_129 br_0_129 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c129
*+ bl_0_129 br_0_129 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c129
*+ bl_0_129 br_0_129 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c129
*+ bl_0_129 br_0_129 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c129
*+ bl_0_129 br_0_129 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c129
*+ bl_0_129 br_0_129 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c129
*+ bl_0_129 br_0_129 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c129
*+ bl_0_129 br_0_129 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c129
*+ bl_0_129 br_0_129 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c129
*+ bl_0_129 br_0_129 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c129
*+ bl_0_129 br_0_129 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c129
*+ bl_0_129 br_0_129 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c129
*+ bl_0_129 br_0_129 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c129
*+ bl_0_129 br_0_129 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c129
*+ bl_0_129 br_0_129 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c129
*+ bl_0_129 br_0_129 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c129
*+ bl_0_129 br_0_129 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c129
*+ bl_0_129 br_0_129 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c129
*+ bl_0_129 br_0_129 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c129
*+ bl_0_129 br_0_129 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c129
+ bl_0_129 br_0_129 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c130
+ bl_0_130 br_0_130 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c130
*+ bl_0_130 br_0_130 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c130
*+ bl_0_130 br_0_130 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c130
*+ bl_0_130 br_0_130 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c130
*+ bl_0_130 br_0_130 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c130
*+ bl_0_130 br_0_130 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c130
*+ bl_0_130 br_0_130 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c130
*+ bl_0_130 br_0_130 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c130
*+ bl_0_130 br_0_130 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c130
*+ bl_0_130 br_0_130 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c130
*+ bl_0_130 br_0_130 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c130
*+ bl_0_130 br_0_130 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c130
*+ bl_0_130 br_0_130 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c130
*+ bl_0_130 br_0_130 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c130
*+ bl_0_130 br_0_130 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c130
*+ bl_0_130 br_0_130 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c130
*+ bl_0_130 br_0_130 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c130
*+ bl_0_130 br_0_130 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c130
*+ bl_0_130 br_0_130 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c130
*+ bl_0_130 br_0_130 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c130
*+ bl_0_130 br_0_130 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c130
*+ bl_0_130 br_0_130 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c130
*+ bl_0_130 br_0_130 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c130
*+ bl_0_130 br_0_130 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c130
*+ bl_0_130 br_0_130 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c130
*+ bl_0_130 br_0_130 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c130
*+ bl_0_130 br_0_130 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c130
*+ bl_0_130 br_0_130 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c130
*+ bl_0_130 br_0_130 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c130
*+ bl_0_130 br_0_130 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c130
*+ bl_0_130 br_0_130 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c130
*+ bl_0_130 br_0_130 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c130
*+ bl_0_130 br_0_130 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c130
*+ bl_0_130 br_0_130 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c130
*+ bl_0_130 br_0_130 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c130
*+ bl_0_130 br_0_130 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c130
*+ bl_0_130 br_0_130 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c130
*+ bl_0_130 br_0_130 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c130
*+ bl_0_130 br_0_130 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c130
*+ bl_0_130 br_0_130 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c130
*+ bl_0_130 br_0_130 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c130
*+ bl_0_130 br_0_130 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c130
*+ bl_0_130 br_0_130 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c130
*+ bl_0_130 br_0_130 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c130
*+ bl_0_130 br_0_130 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c130
*+ bl_0_130 br_0_130 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c130
*+ bl_0_130 br_0_130 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c130
*+ bl_0_130 br_0_130 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c130
*+ bl_0_130 br_0_130 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c130
*+ bl_0_130 br_0_130 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c130
*+ bl_0_130 br_0_130 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c130
*+ bl_0_130 br_0_130 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c130
*+ bl_0_130 br_0_130 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c130
*+ bl_0_130 br_0_130 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c130
*+ bl_0_130 br_0_130 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c130
*+ bl_0_130 br_0_130 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c130
*+ bl_0_130 br_0_130 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c130
*+ bl_0_130 br_0_130 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c130
*+ bl_0_130 br_0_130 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c130
*+ bl_0_130 br_0_130 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c130
*+ bl_0_130 br_0_130 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c130
*+ bl_0_130 br_0_130 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c130
*+ bl_0_130 br_0_130 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c130
*+ bl_0_130 br_0_130 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c130
*+ bl_0_130 br_0_130 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c130
*+ bl_0_130 br_0_130 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c130
*+ bl_0_130 br_0_130 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c130
*+ bl_0_130 br_0_130 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c130
*+ bl_0_130 br_0_130 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c130
*+ bl_0_130 br_0_130 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c130
*+ bl_0_130 br_0_130 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c130
*+ bl_0_130 br_0_130 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c130
*+ bl_0_130 br_0_130 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c130
*+ bl_0_130 br_0_130 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c130
*+ bl_0_130 br_0_130 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c130
*+ bl_0_130 br_0_130 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c130
*+ bl_0_130 br_0_130 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c130
*+ bl_0_130 br_0_130 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c130
*+ bl_0_130 br_0_130 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c130
*+ bl_0_130 br_0_130 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c130
*+ bl_0_130 br_0_130 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c130
*+ bl_0_130 br_0_130 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c130
*+ bl_0_130 br_0_130 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c130
*+ bl_0_130 br_0_130 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c130
*+ bl_0_130 br_0_130 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c130
*+ bl_0_130 br_0_130 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c130
*+ bl_0_130 br_0_130 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c130
*+ bl_0_130 br_0_130 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c130
*+ bl_0_130 br_0_130 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c130
*+ bl_0_130 br_0_130 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c130
*+ bl_0_130 br_0_130 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c130
*+ bl_0_130 br_0_130 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c130
*+ bl_0_130 br_0_130 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c130
*+ bl_0_130 br_0_130 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c130
*+ bl_0_130 br_0_130 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c130
*+ bl_0_130 br_0_130 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c130
*+ bl_0_130 br_0_130 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c130
*+ bl_0_130 br_0_130 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c130
*+ bl_0_130 br_0_130 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c130
*+ bl_0_130 br_0_130 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c130
*+ bl_0_130 br_0_130 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c130
*+ bl_0_130 br_0_130 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c130
*+ bl_0_130 br_0_130 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c130
*+ bl_0_130 br_0_130 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c130
*+ bl_0_130 br_0_130 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c130
*+ bl_0_130 br_0_130 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c130
*+ bl_0_130 br_0_130 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c130
*+ bl_0_130 br_0_130 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c130
*+ bl_0_130 br_0_130 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c130
*+ bl_0_130 br_0_130 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c130
*+ bl_0_130 br_0_130 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c130
*+ bl_0_130 br_0_130 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c130
*+ bl_0_130 br_0_130 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c130
*+ bl_0_130 br_0_130 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c130
*+ bl_0_130 br_0_130 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c130
*+ bl_0_130 br_0_130 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c130
*+ bl_0_130 br_0_130 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c130
*+ bl_0_130 br_0_130 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c130
*+ bl_0_130 br_0_130 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c130
*+ bl_0_130 br_0_130 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c130
*+ bl_0_130 br_0_130 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c130
*+ bl_0_130 br_0_130 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c130
*+ bl_0_130 br_0_130 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c130
*+ bl_0_130 br_0_130 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c130
*+ bl_0_130 br_0_130 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c130
*+ bl_0_130 br_0_130 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c130
*+ bl_0_130 br_0_130 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c130
+ bl_0_130 br_0_130 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c131
+ bl_0_131 br_0_131 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c131
*+ bl_0_131 br_0_131 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c131
*+ bl_0_131 br_0_131 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c131
*+ bl_0_131 br_0_131 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c131
*+ bl_0_131 br_0_131 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c131
*+ bl_0_131 br_0_131 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c131
*+ bl_0_131 br_0_131 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c131
*+ bl_0_131 br_0_131 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c131
*+ bl_0_131 br_0_131 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c131
*+ bl_0_131 br_0_131 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c131
*+ bl_0_131 br_0_131 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c131
*+ bl_0_131 br_0_131 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c131
*+ bl_0_131 br_0_131 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c131
*+ bl_0_131 br_0_131 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c131
*+ bl_0_131 br_0_131 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c131
*+ bl_0_131 br_0_131 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c131
*+ bl_0_131 br_0_131 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c131
*+ bl_0_131 br_0_131 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c131
*+ bl_0_131 br_0_131 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c131
*+ bl_0_131 br_0_131 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c131
*+ bl_0_131 br_0_131 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c131
*+ bl_0_131 br_0_131 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c131
*+ bl_0_131 br_0_131 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c131
*+ bl_0_131 br_0_131 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c131
*+ bl_0_131 br_0_131 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c131
*+ bl_0_131 br_0_131 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c131
*+ bl_0_131 br_0_131 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c131
*+ bl_0_131 br_0_131 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c131
*+ bl_0_131 br_0_131 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c131
*+ bl_0_131 br_0_131 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c131
*+ bl_0_131 br_0_131 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c131
*+ bl_0_131 br_0_131 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c131
*+ bl_0_131 br_0_131 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c131
*+ bl_0_131 br_0_131 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c131
*+ bl_0_131 br_0_131 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c131
*+ bl_0_131 br_0_131 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c131
*+ bl_0_131 br_0_131 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c131
*+ bl_0_131 br_0_131 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c131
*+ bl_0_131 br_0_131 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c131
*+ bl_0_131 br_0_131 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c131
*+ bl_0_131 br_0_131 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c131
*+ bl_0_131 br_0_131 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c131
*+ bl_0_131 br_0_131 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c131
*+ bl_0_131 br_0_131 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c131
*+ bl_0_131 br_0_131 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c131
*+ bl_0_131 br_0_131 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c131
*+ bl_0_131 br_0_131 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c131
*+ bl_0_131 br_0_131 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c131
*+ bl_0_131 br_0_131 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c131
*+ bl_0_131 br_0_131 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c131
*+ bl_0_131 br_0_131 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c131
*+ bl_0_131 br_0_131 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c131
*+ bl_0_131 br_0_131 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c131
*+ bl_0_131 br_0_131 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c131
*+ bl_0_131 br_0_131 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c131
*+ bl_0_131 br_0_131 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c131
*+ bl_0_131 br_0_131 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c131
*+ bl_0_131 br_0_131 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c131
*+ bl_0_131 br_0_131 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c131
*+ bl_0_131 br_0_131 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c131
*+ bl_0_131 br_0_131 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c131
*+ bl_0_131 br_0_131 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c131
*+ bl_0_131 br_0_131 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c131
*+ bl_0_131 br_0_131 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c131
*+ bl_0_131 br_0_131 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c131
*+ bl_0_131 br_0_131 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c131
*+ bl_0_131 br_0_131 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c131
*+ bl_0_131 br_0_131 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c131
*+ bl_0_131 br_0_131 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c131
*+ bl_0_131 br_0_131 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c131
*+ bl_0_131 br_0_131 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c131
*+ bl_0_131 br_0_131 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c131
*+ bl_0_131 br_0_131 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c131
*+ bl_0_131 br_0_131 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c131
*+ bl_0_131 br_0_131 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c131
*+ bl_0_131 br_0_131 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c131
*+ bl_0_131 br_0_131 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c131
*+ bl_0_131 br_0_131 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c131
*+ bl_0_131 br_0_131 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c131
*+ bl_0_131 br_0_131 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c131
*+ bl_0_131 br_0_131 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c131
*+ bl_0_131 br_0_131 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c131
*+ bl_0_131 br_0_131 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c131
*+ bl_0_131 br_0_131 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c131
*+ bl_0_131 br_0_131 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c131
*+ bl_0_131 br_0_131 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c131
*+ bl_0_131 br_0_131 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c131
*+ bl_0_131 br_0_131 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c131
*+ bl_0_131 br_0_131 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c131
*+ bl_0_131 br_0_131 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c131
*+ bl_0_131 br_0_131 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c131
*+ bl_0_131 br_0_131 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c131
*+ bl_0_131 br_0_131 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c131
*+ bl_0_131 br_0_131 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c131
*+ bl_0_131 br_0_131 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c131
*+ bl_0_131 br_0_131 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c131
*+ bl_0_131 br_0_131 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c131
*+ bl_0_131 br_0_131 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c131
*+ bl_0_131 br_0_131 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c131
*+ bl_0_131 br_0_131 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c131
*+ bl_0_131 br_0_131 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c131
*+ bl_0_131 br_0_131 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c131
*+ bl_0_131 br_0_131 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c131
*+ bl_0_131 br_0_131 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c131
*+ bl_0_131 br_0_131 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c131
*+ bl_0_131 br_0_131 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c131
*+ bl_0_131 br_0_131 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c131
*+ bl_0_131 br_0_131 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c131
*+ bl_0_131 br_0_131 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c131
*+ bl_0_131 br_0_131 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c131
*+ bl_0_131 br_0_131 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c131
*+ bl_0_131 br_0_131 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c131
*+ bl_0_131 br_0_131 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c131
*+ bl_0_131 br_0_131 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c131
*+ bl_0_131 br_0_131 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c131
*+ bl_0_131 br_0_131 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c131
*+ bl_0_131 br_0_131 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c131
*+ bl_0_131 br_0_131 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c131
*+ bl_0_131 br_0_131 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c131
*+ bl_0_131 br_0_131 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c131
*+ bl_0_131 br_0_131 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c131
*+ bl_0_131 br_0_131 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c131
*+ bl_0_131 br_0_131 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c131
*+ bl_0_131 br_0_131 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c131
*+ bl_0_131 br_0_131 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c131
*+ bl_0_131 br_0_131 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c131
*+ bl_0_131 br_0_131 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c131
+ bl_0_131 br_0_131 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c132
+ bl_0_132 br_0_132 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c132
*+ bl_0_132 br_0_132 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c132
*+ bl_0_132 br_0_132 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c132
*+ bl_0_132 br_0_132 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c132
*+ bl_0_132 br_0_132 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c132
*+ bl_0_132 br_0_132 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c132
*+ bl_0_132 br_0_132 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c132
*+ bl_0_132 br_0_132 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c132
*+ bl_0_132 br_0_132 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c132
*+ bl_0_132 br_0_132 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c132
*+ bl_0_132 br_0_132 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c132
*+ bl_0_132 br_0_132 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c132
*+ bl_0_132 br_0_132 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c132
*+ bl_0_132 br_0_132 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c132
*+ bl_0_132 br_0_132 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c132
*+ bl_0_132 br_0_132 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c132
*+ bl_0_132 br_0_132 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c132
*+ bl_0_132 br_0_132 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c132
*+ bl_0_132 br_0_132 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c132
*+ bl_0_132 br_0_132 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c132
*+ bl_0_132 br_0_132 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c132
*+ bl_0_132 br_0_132 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c132
*+ bl_0_132 br_0_132 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c132
*+ bl_0_132 br_0_132 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c132
*+ bl_0_132 br_0_132 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c132
*+ bl_0_132 br_0_132 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c132
*+ bl_0_132 br_0_132 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c132
*+ bl_0_132 br_0_132 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c132
*+ bl_0_132 br_0_132 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c132
*+ bl_0_132 br_0_132 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c132
*+ bl_0_132 br_0_132 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c132
*+ bl_0_132 br_0_132 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c132
*+ bl_0_132 br_0_132 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c132
*+ bl_0_132 br_0_132 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c132
*+ bl_0_132 br_0_132 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c132
*+ bl_0_132 br_0_132 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c132
*+ bl_0_132 br_0_132 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c132
*+ bl_0_132 br_0_132 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c132
*+ bl_0_132 br_0_132 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c132
*+ bl_0_132 br_0_132 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c132
*+ bl_0_132 br_0_132 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c132
*+ bl_0_132 br_0_132 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c132
*+ bl_0_132 br_0_132 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c132
*+ bl_0_132 br_0_132 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c132
*+ bl_0_132 br_0_132 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c132
*+ bl_0_132 br_0_132 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c132
*+ bl_0_132 br_0_132 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c132
*+ bl_0_132 br_0_132 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c132
*+ bl_0_132 br_0_132 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c132
*+ bl_0_132 br_0_132 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c132
*+ bl_0_132 br_0_132 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c132
*+ bl_0_132 br_0_132 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c132
*+ bl_0_132 br_0_132 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c132
*+ bl_0_132 br_0_132 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c132
*+ bl_0_132 br_0_132 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c132
*+ bl_0_132 br_0_132 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c132
*+ bl_0_132 br_0_132 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c132
*+ bl_0_132 br_0_132 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c132
*+ bl_0_132 br_0_132 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c132
*+ bl_0_132 br_0_132 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c132
*+ bl_0_132 br_0_132 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c132
*+ bl_0_132 br_0_132 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c132
*+ bl_0_132 br_0_132 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c132
*+ bl_0_132 br_0_132 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c132
*+ bl_0_132 br_0_132 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c132
*+ bl_0_132 br_0_132 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c132
*+ bl_0_132 br_0_132 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c132
*+ bl_0_132 br_0_132 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c132
*+ bl_0_132 br_0_132 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c132
*+ bl_0_132 br_0_132 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c132
*+ bl_0_132 br_0_132 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c132
*+ bl_0_132 br_0_132 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c132
*+ bl_0_132 br_0_132 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c132
*+ bl_0_132 br_0_132 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c132
*+ bl_0_132 br_0_132 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c132
*+ bl_0_132 br_0_132 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c132
*+ bl_0_132 br_0_132 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c132
*+ bl_0_132 br_0_132 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c132
*+ bl_0_132 br_0_132 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c132
*+ bl_0_132 br_0_132 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c132
*+ bl_0_132 br_0_132 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c132
*+ bl_0_132 br_0_132 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c132
*+ bl_0_132 br_0_132 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c132
*+ bl_0_132 br_0_132 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c132
*+ bl_0_132 br_0_132 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c132
*+ bl_0_132 br_0_132 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c132
*+ bl_0_132 br_0_132 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c132
*+ bl_0_132 br_0_132 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c132
*+ bl_0_132 br_0_132 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c132
*+ bl_0_132 br_0_132 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c132
*+ bl_0_132 br_0_132 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c132
*+ bl_0_132 br_0_132 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c132
*+ bl_0_132 br_0_132 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c132
*+ bl_0_132 br_0_132 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c132
*+ bl_0_132 br_0_132 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c132
*+ bl_0_132 br_0_132 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c132
*+ bl_0_132 br_0_132 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c132
*+ bl_0_132 br_0_132 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c132
*+ bl_0_132 br_0_132 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c132
*+ bl_0_132 br_0_132 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c132
*+ bl_0_132 br_0_132 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c132
*+ bl_0_132 br_0_132 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c132
*+ bl_0_132 br_0_132 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c132
*+ bl_0_132 br_0_132 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c132
*+ bl_0_132 br_0_132 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c132
*+ bl_0_132 br_0_132 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c132
*+ bl_0_132 br_0_132 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c132
*+ bl_0_132 br_0_132 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c132
*+ bl_0_132 br_0_132 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c132
*+ bl_0_132 br_0_132 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c132
*+ bl_0_132 br_0_132 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c132
*+ bl_0_132 br_0_132 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c132
*+ bl_0_132 br_0_132 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c132
*+ bl_0_132 br_0_132 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c132
*+ bl_0_132 br_0_132 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c132
*+ bl_0_132 br_0_132 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c132
*+ bl_0_132 br_0_132 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c132
*+ bl_0_132 br_0_132 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c132
*+ bl_0_132 br_0_132 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c132
*+ bl_0_132 br_0_132 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c132
*+ bl_0_132 br_0_132 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c132
*+ bl_0_132 br_0_132 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c132
*+ bl_0_132 br_0_132 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c132
*+ bl_0_132 br_0_132 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c132
*+ bl_0_132 br_0_132 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c132
*+ bl_0_132 br_0_132 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c132
*+ bl_0_132 br_0_132 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c132
+ bl_0_132 br_0_132 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c133
+ bl_0_133 br_0_133 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c133
*+ bl_0_133 br_0_133 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c133
*+ bl_0_133 br_0_133 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c133
*+ bl_0_133 br_0_133 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c133
*+ bl_0_133 br_0_133 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c133
*+ bl_0_133 br_0_133 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c133
*+ bl_0_133 br_0_133 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c133
*+ bl_0_133 br_0_133 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c133
*+ bl_0_133 br_0_133 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c133
*+ bl_0_133 br_0_133 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c133
*+ bl_0_133 br_0_133 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c133
*+ bl_0_133 br_0_133 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c133
*+ bl_0_133 br_0_133 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c133
*+ bl_0_133 br_0_133 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c133
*+ bl_0_133 br_0_133 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c133
*+ bl_0_133 br_0_133 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c133
*+ bl_0_133 br_0_133 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c133
*+ bl_0_133 br_0_133 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c133
*+ bl_0_133 br_0_133 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c133
*+ bl_0_133 br_0_133 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c133
*+ bl_0_133 br_0_133 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c133
*+ bl_0_133 br_0_133 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c133
*+ bl_0_133 br_0_133 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c133
*+ bl_0_133 br_0_133 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c133
*+ bl_0_133 br_0_133 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c133
*+ bl_0_133 br_0_133 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c133
*+ bl_0_133 br_0_133 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c133
*+ bl_0_133 br_0_133 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c133
*+ bl_0_133 br_0_133 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c133
*+ bl_0_133 br_0_133 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c133
*+ bl_0_133 br_0_133 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c133
*+ bl_0_133 br_0_133 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c133
*+ bl_0_133 br_0_133 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c133
*+ bl_0_133 br_0_133 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c133
*+ bl_0_133 br_0_133 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c133
*+ bl_0_133 br_0_133 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c133
*+ bl_0_133 br_0_133 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c133
*+ bl_0_133 br_0_133 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c133
*+ bl_0_133 br_0_133 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c133
*+ bl_0_133 br_0_133 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c133
*+ bl_0_133 br_0_133 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c133
*+ bl_0_133 br_0_133 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c133
*+ bl_0_133 br_0_133 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c133
*+ bl_0_133 br_0_133 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c133
*+ bl_0_133 br_0_133 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c133
*+ bl_0_133 br_0_133 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c133
*+ bl_0_133 br_0_133 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c133
*+ bl_0_133 br_0_133 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c133
*+ bl_0_133 br_0_133 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c133
*+ bl_0_133 br_0_133 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c133
*+ bl_0_133 br_0_133 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c133
*+ bl_0_133 br_0_133 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c133
*+ bl_0_133 br_0_133 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c133
*+ bl_0_133 br_0_133 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c133
*+ bl_0_133 br_0_133 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c133
*+ bl_0_133 br_0_133 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c133
*+ bl_0_133 br_0_133 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c133
*+ bl_0_133 br_0_133 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c133
*+ bl_0_133 br_0_133 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c133
*+ bl_0_133 br_0_133 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c133
*+ bl_0_133 br_0_133 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c133
*+ bl_0_133 br_0_133 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c133
*+ bl_0_133 br_0_133 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c133
*+ bl_0_133 br_0_133 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c133
*+ bl_0_133 br_0_133 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c133
*+ bl_0_133 br_0_133 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c133
*+ bl_0_133 br_0_133 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c133
*+ bl_0_133 br_0_133 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c133
*+ bl_0_133 br_0_133 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c133
*+ bl_0_133 br_0_133 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c133
*+ bl_0_133 br_0_133 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c133
*+ bl_0_133 br_0_133 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c133
*+ bl_0_133 br_0_133 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c133
*+ bl_0_133 br_0_133 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c133
*+ bl_0_133 br_0_133 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c133
*+ bl_0_133 br_0_133 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c133
*+ bl_0_133 br_0_133 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c133
*+ bl_0_133 br_0_133 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c133
*+ bl_0_133 br_0_133 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c133
*+ bl_0_133 br_0_133 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c133
*+ bl_0_133 br_0_133 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c133
*+ bl_0_133 br_0_133 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c133
*+ bl_0_133 br_0_133 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c133
*+ bl_0_133 br_0_133 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c133
*+ bl_0_133 br_0_133 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c133
*+ bl_0_133 br_0_133 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c133
*+ bl_0_133 br_0_133 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c133
*+ bl_0_133 br_0_133 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c133
*+ bl_0_133 br_0_133 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c133
*+ bl_0_133 br_0_133 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c133
*+ bl_0_133 br_0_133 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c133
*+ bl_0_133 br_0_133 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c133
*+ bl_0_133 br_0_133 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c133
*+ bl_0_133 br_0_133 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c133
*+ bl_0_133 br_0_133 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c133
*+ bl_0_133 br_0_133 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c133
*+ bl_0_133 br_0_133 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c133
*+ bl_0_133 br_0_133 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c133
*+ bl_0_133 br_0_133 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c133
*+ bl_0_133 br_0_133 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c133
*+ bl_0_133 br_0_133 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c133
*+ bl_0_133 br_0_133 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c133
*+ bl_0_133 br_0_133 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c133
*+ bl_0_133 br_0_133 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c133
*+ bl_0_133 br_0_133 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c133
*+ bl_0_133 br_0_133 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c133
*+ bl_0_133 br_0_133 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c133
*+ bl_0_133 br_0_133 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c133
*+ bl_0_133 br_0_133 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c133
*+ bl_0_133 br_0_133 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c133
*+ bl_0_133 br_0_133 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c133
*+ bl_0_133 br_0_133 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c133
*+ bl_0_133 br_0_133 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c133
*+ bl_0_133 br_0_133 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c133
*+ bl_0_133 br_0_133 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c133
*+ bl_0_133 br_0_133 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c133
*+ bl_0_133 br_0_133 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c133
*+ bl_0_133 br_0_133 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c133
*+ bl_0_133 br_0_133 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c133
*+ bl_0_133 br_0_133 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c133
*+ bl_0_133 br_0_133 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c133
*+ bl_0_133 br_0_133 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c133
*+ bl_0_133 br_0_133 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c133
*+ bl_0_133 br_0_133 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c133
*+ bl_0_133 br_0_133 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c133
*+ bl_0_133 br_0_133 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c133
*+ bl_0_133 br_0_133 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c133
+ bl_0_133 br_0_133 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c134
+ bl_0_134 br_0_134 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c134
*+ bl_0_134 br_0_134 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c134
*+ bl_0_134 br_0_134 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c134
*+ bl_0_134 br_0_134 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c134
*+ bl_0_134 br_0_134 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c134
*+ bl_0_134 br_0_134 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c134
*+ bl_0_134 br_0_134 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c134
*+ bl_0_134 br_0_134 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c134
*+ bl_0_134 br_0_134 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c134
*+ bl_0_134 br_0_134 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c134
*+ bl_0_134 br_0_134 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c134
*+ bl_0_134 br_0_134 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c134
*+ bl_0_134 br_0_134 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c134
*+ bl_0_134 br_0_134 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c134
*+ bl_0_134 br_0_134 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c134
*+ bl_0_134 br_0_134 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c134
*+ bl_0_134 br_0_134 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c134
*+ bl_0_134 br_0_134 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c134
*+ bl_0_134 br_0_134 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c134
*+ bl_0_134 br_0_134 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c134
*+ bl_0_134 br_0_134 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c134
*+ bl_0_134 br_0_134 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c134
*+ bl_0_134 br_0_134 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c134
*+ bl_0_134 br_0_134 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c134
*+ bl_0_134 br_0_134 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c134
*+ bl_0_134 br_0_134 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c134
*+ bl_0_134 br_0_134 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c134
*+ bl_0_134 br_0_134 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c134
*+ bl_0_134 br_0_134 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c134
*+ bl_0_134 br_0_134 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c134
*+ bl_0_134 br_0_134 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c134
*+ bl_0_134 br_0_134 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c134
*+ bl_0_134 br_0_134 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c134
*+ bl_0_134 br_0_134 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c134
*+ bl_0_134 br_0_134 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c134
*+ bl_0_134 br_0_134 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c134
*+ bl_0_134 br_0_134 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c134
*+ bl_0_134 br_0_134 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c134
*+ bl_0_134 br_0_134 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c134
*+ bl_0_134 br_0_134 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c134
*+ bl_0_134 br_0_134 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c134
*+ bl_0_134 br_0_134 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c134
*+ bl_0_134 br_0_134 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c134
*+ bl_0_134 br_0_134 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c134
*+ bl_0_134 br_0_134 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c134
*+ bl_0_134 br_0_134 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c134
*+ bl_0_134 br_0_134 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c134
*+ bl_0_134 br_0_134 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c134
*+ bl_0_134 br_0_134 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c134
*+ bl_0_134 br_0_134 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c134
*+ bl_0_134 br_0_134 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c134
*+ bl_0_134 br_0_134 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c134
*+ bl_0_134 br_0_134 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c134
*+ bl_0_134 br_0_134 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c134
*+ bl_0_134 br_0_134 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c134
*+ bl_0_134 br_0_134 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c134
*+ bl_0_134 br_0_134 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c134
*+ bl_0_134 br_0_134 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c134
*+ bl_0_134 br_0_134 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c134
*+ bl_0_134 br_0_134 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c134
*+ bl_0_134 br_0_134 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c134
*+ bl_0_134 br_0_134 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c134
*+ bl_0_134 br_0_134 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c134
*+ bl_0_134 br_0_134 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c134
*+ bl_0_134 br_0_134 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c134
*+ bl_0_134 br_0_134 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c134
*+ bl_0_134 br_0_134 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c134
*+ bl_0_134 br_0_134 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c134
*+ bl_0_134 br_0_134 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c134
*+ bl_0_134 br_0_134 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c134
*+ bl_0_134 br_0_134 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c134
*+ bl_0_134 br_0_134 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c134
*+ bl_0_134 br_0_134 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c134
*+ bl_0_134 br_0_134 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c134
*+ bl_0_134 br_0_134 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c134
*+ bl_0_134 br_0_134 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c134
*+ bl_0_134 br_0_134 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c134
*+ bl_0_134 br_0_134 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c134
*+ bl_0_134 br_0_134 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c134
*+ bl_0_134 br_0_134 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c134
*+ bl_0_134 br_0_134 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c134
*+ bl_0_134 br_0_134 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c134
*+ bl_0_134 br_0_134 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c134
*+ bl_0_134 br_0_134 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c134
*+ bl_0_134 br_0_134 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c134
*+ bl_0_134 br_0_134 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c134
*+ bl_0_134 br_0_134 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c134
*+ bl_0_134 br_0_134 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c134
*+ bl_0_134 br_0_134 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c134
*+ bl_0_134 br_0_134 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c134
*+ bl_0_134 br_0_134 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c134
*+ bl_0_134 br_0_134 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c134
*+ bl_0_134 br_0_134 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c134
*+ bl_0_134 br_0_134 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c134
*+ bl_0_134 br_0_134 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c134
*+ bl_0_134 br_0_134 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c134
*+ bl_0_134 br_0_134 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c134
*+ bl_0_134 br_0_134 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c134
*+ bl_0_134 br_0_134 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c134
*+ bl_0_134 br_0_134 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c134
*+ bl_0_134 br_0_134 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c134
*+ bl_0_134 br_0_134 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c134
*+ bl_0_134 br_0_134 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c134
*+ bl_0_134 br_0_134 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c134
*+ bl_0_134 br_0_134 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c134
*+ bl_0_134 br_0_134 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c134
*+ bl_0_134 br_0_134 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c134
*+ bl_0_134 br_0_134 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c134
*+ bl_0_134 br_0_134 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c134
*+ bl_0_134 br_0_134 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c134
*+ bl_0_134 br_0_134 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c134
*+ bl_0_134 br_0_134 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c134
*+ bl_0_134 br_0_134 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c134
*+ bl_0_134 br_0_134 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c134
*+ bl_0_134 br_0_134 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c134
*+ bl_0_134 br_0_134 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c134
*+ bl_0_134 br_0_134 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c134
*+ bl_0_134 br_0_134 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c134
*+ bl_0_134 br_0_134 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c134
*+ bl_0_134 br_0_134 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c134
*+ bl_0_134 br_0_134 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c134
*+ bl_0_134 br_0_134 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c134
*+ bl_0_134 br_0_134 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c134
*+ bl_0_134 br_0_134 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c134
*+ bl_0_134 br_0_134 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c134
*+ bl_0_134 br_0_134 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c134
*+ bl_0_134 br_0_134 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c134
+ bl_0_134 br_0_134 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c135
+ bl_0_135 br_0_135 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c135
*+ bl_0_135 br_0_135 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c135
*+ bl_0_135 br_0_135 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c135
*+ bl_0_135 br_0_135 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c135
*+ bl_0_135 br_0_135 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c135
*+ bl_0_135 br_0_135 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c135
*+ bl_0_135 br_0_135 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c135
*+ bl_0_135 br_0_135 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c135
*+ bl_0_135 br_0_135 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c135
*+ bl_0_135 br_0_135 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c135
*+ bl_0_135 br_0_135 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c135
*+ bl_0_135 br_0_135 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c135
*+ bl_0_135 br_0_135 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c135
*+ bl_0_135 br_0_135 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c135
*+ bl_0_135 br_0_135 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c135
*+ bl_0_135 br_0_135 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c135
*+ bl_0_135 br_0_135 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c135
*+ bl_0_135 br_0_135 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c135
*+ bl_0_135 br_0_135 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c135
*+ bl_0_135 br_0_135 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c135
*+ bl_0_135 br_0_135 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c135
*+ bl_0_135 br_0_135 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c135
*+ bl_0_135 br_0_135 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c135
*+ bl_0_135 br_0_135 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c135
*+ bl_0_135 br_0_135 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c135
*+ bl_0_135 br_0_135 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c135
*+ bl_0_135 br_0_135 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c135
*+ bl_0_135 br_0_135 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c135
*+ bl_0_135 br_0_135 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c135
*+ bl_0_135 br_0_135 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c135
*+ bl_0_135 br_0_135 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c135
*+ bl_0_135 br_0_135 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c135
*+ bl_0_135 br_0_135 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c135
*+ bl_0_135 br_0_135 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c135
*+ bl_0_135 br_0_135 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c135
*+ bl_0_135 br_0_135 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c135
*+ bl_0_135 br_0_135 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c135
*+ bl_0_135 br_0_135 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c135
*+ bl_0_135 br_0_135 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c135
*+ bl_0_135 br_0_135 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c135
*+ bl_0_135 br_0_135 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c135
*+ bl_0_135 br_0_135 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c135
*+ bl_0_135 br_0_135 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c135
*+ bl_0_135 br_0_135 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c135
*+ bl_0_135 br_0_135 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c135
*+ bl_0_135 br_0_135 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c135
*+ bl_0_135 br_0_135 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c135
*+ bl_0_135 br_0_135 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c135
*+ bl_0_135 br_0_135 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c135
*+ bl_0_135 br_0_135 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c135
*+ bl_0_135 br_0_135 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c135
*+ bl_0_135 br_0_135 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c135
*+ bl_0_135 br_0_135 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c135
*+ bl_0_135 br_0_135 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c135
*+ bl_0_135 br_0_135 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c135
*+ bl_0_135 br_0_135 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c135
*+ bl_0_135 br_0_135 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c135
*+ bl_0_135 br_0_135 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c135
*+ bl_0_135 br_0_135 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c135
*+ bl_0_135 br_0_135 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c135
*+ bl_0_135 br_0_135 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c135
*+ bl_0_135 br_0_135 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c135
*+ bl_0_135 br_0_135 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c135
*+ bl_0_135 br_0_135 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c135
*+ bl_0_135 br_0_135 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c135
*+ bl_0_135 br_0_135 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c135
*+ bl_0_135 br_0_135 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c135
*+ bl_0_135 br_0_135 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c135
*+ bl_0_135 br_0_135 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c135
*+ bl_0_135 br_0_135 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c135
*+ bl_0_135 br_0_135 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c135
*+ bl_0_135 br_0_135 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c135
*+ bl_0_135 br_0_135 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c135
*+ bl_0_135 br_0_135 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c135
*+ bl_0_135 br_0_135 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c135
*+ bl_0_135 br_0_135 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c135
*+ bl_0_135 br_0_135 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c135
*+ bl_0_135 br_0_135 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c135
*+ bl_0_135 br_0_135 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c135
*+ bl_0_135 br_0_135 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c135
*+ bl_0_135 br_0_135 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c135
*+ bl_0_135 br_0_135 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c135
*+ bl_0_135 br_0_135 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c135
*+ bl_0_135 br_0_135 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c135
*+ bl_0_135 br_0_135 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c135
*+ bl_0_135 br_0_135 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c135
*+ bl_0_135 br_0_135 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c135
*+ bl_0_135 br_0_135 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c135
*+ bl_0_135 br_0_135 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c135
*+ bl_0_135 br_0_135 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c135
*+ bl_0_135 br_0_135 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c135
*+ bl_0_135 br_0_135 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c135
*+ bl_0_135 br_0_135 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c135
*+ bl_0_135 br_0_135 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c135
*+ bl_0_135 br_0_135 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c135
*+ bl_0_135 br_0_135 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c135
*+ bl_0_135 br_0_135 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c135
*+ bl_0_135 br_0_135 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c135
*+ bl_0_135 br_0_135 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c135
*+ bl_0_135 br_0_135 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c135
*+ bl_0_135 br_0_135 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c135
*+ bl_0_135 br_0_135 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c135
*+ bl_0_135 br_0_135 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c135
*+ bl_0_135 br_0_135 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c135
*+ bl_0_135 br_0_135 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c135
*+ bl_0_135 br_0_135 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c135
*+ bl_0_135 br_0_135 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c135
*+ bl_0_135 br_0_135 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c135
*+ bl_0_135 br_0_135 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c135
*+ bl_0_135 br_0_135 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c135
*+ bl_0_135 br_0_135 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c135
*+ bl_0_135 br_0_135 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c135
*+ bl_0_135 br_0_135 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c135
*+ bl_0_135 br_0_135 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c135
*+ bl_0_135 br_0_135 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c135
*+ bl_0_135 br_0_135 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c135
*+ bl_0_135 br_0_135 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c135
*+ bl_0_135 br_0_135 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c135
*+ bl_0_135 br_0_135 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c135
*+ bl_0_135 br_0_135 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c135
*+ bl_0_135 br_0_135 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c135
*+ bl_0_135 br_0_135 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c135
*+ bl_0_135 br_0_135 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c135
*+ bl_0_135 br_0_135 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c135
*+ bl_0_135 br_0_135 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c135
*+ bl_0_135 br_0_135 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c135
*+ bl_0_135 br_0_135 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c135
+ bl_0_135 br_0_135 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c136
+ bl_0_136 br_0_136 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c136
*+ bl_0_136 br_0_136 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c136
*+ bl_0_136 br_0_136 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c136
*+ bl_0_136 br_0_136 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c136
*+ bl_0_136 br_0_136 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c136
*+ bl_0_136 br_0_136 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c136
*+ bl_0_136 br_0_136 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c136
*+ bl_0_136 br_0_136 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c136
*+ bl_0_136 br_0_136 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c136
*+ bl_0_136 br_0_136 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c136
*+ bl_0_136 br_0_136 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c136
*+ bl_0_136 br_0_136 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c136
*+ bl_0_136 br_0_136 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c136
*+ bl_0_136 br_0_136 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c136
*+ bl_0_136 br_0_136 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c136
*+ bl_0_136 br_0_136 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c136
*+ bl_0_136 br_0_136 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c136
*+ bl_0_136 br_0_136 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c136
*+ bl_0_136 br_0_136 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c136
*+ bl_0_136 br_0_136 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c136
*+ bl_0_136 br_0_136 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c136
*+ bl_0_136 br_0_136 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c136
*+ bl_0_136 br_0_136 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c136
*+ bl_0_136 br_0_136 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c136
*+ bl_0_136 br_0_136 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c136
*+ bl_0_136 br_0_136 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c136
*+ bl_0_136 br_0_136 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c136
*+ bl_0_136 br_0_136 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c136
*+ bl_0_136 br_0_136 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c136
*+ bl_0_136 br_0_136 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c136
*+ bl_0_136 br_0_136 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c136
*+ bl_0_136 br_0_136 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c136
*+ bl_0_136 br_0_136 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c136
*+ bl_0_136 br_0_136 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c136
*+ bl_0_136 br_0_136 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c136
*+ bl_0_136 br_0_136 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c136
*+ bl_0_136 br_0_136 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c136
*+ bl_0_136 br_0_136 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c136
*+ bl_0_136 br_0_136 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c136
*+ bl_0_136 br_0_136 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c136
*+ bl_0_136 br_0_136 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c136
*+ bl_0_136 br_0_136 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c136
*+ bl_0_136 br_0_136 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c136
*+ bl_0_136 br_0_136 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c136
*+ bl_0_136 br_0_136 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c136
*+ bl_0_136 br_0_136 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c136
*+ bl_0_136 br_0_136 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c136
*+ bl_0_136 br_0_136 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c136
*+ bl_0_136 br_0_136 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c136
*+ bl_0_136 br_0_136 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c136
*+ bl_0_136 br_0_136 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c136
*+ bl_0_136 br_0_136 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c136
*+ bl_0_136 br_0_136 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c136
*+ bl_0_136 br_0_136 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c136
*+ bl_0_136 br_0_136 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c136
*+ bl_0_136 br_0_136 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c136
*+ bl_0_136 br_0_136 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c136
*+ bl_0_136 br_0_136 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c136
*+ bl_0_136 br_0_136 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c136
*+ bl_0_136 br_0_136 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c136
*+ bl_0_136 br_0_136 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c136
*+ bl_0_136 br_0_136 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c136
*+ bl_0_136 br_0_136 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c136
*+ bl_0_136 br_0_136 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c136
*+ bl_0_136 br_0_136 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c136
*+ bl_0_136 br_0_136 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c136
*+ bl_0_136 br_0_136 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c136
*+ bl_0_136 br_0_136 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c136
*+ bl_0_136 br_0_136 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c136
*+ bl_0_136 br_0_136 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c136
*+ bl_0_136 br_0_136 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c136
*+ bl_0_136 br_0_136 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c136
*+ bl_0_136 br_0_136 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c136
*+ bl_0_136 br_0_136 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c136
*+ bl_0_136 br_0_136 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c136
*+ bl_0_136 br_0_136 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c136
*+ bl_0_136 br_0_136 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c136
*+ bl_0_136 br_0_136 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c136
*+ bl_0_136 br_0_136 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c136
*+ bl_0_136 br_0_136 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c136
*+ bl_0_136 br_0_136 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c136
*+ bl_0_136 br_0_136 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c136
*+ bl_0_136 br_0_136 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c136
*+ bl_0_136 br_0_136 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c136
*+ bl_0_136 br_0_136 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c136
*+ bl_0_136 br_0_136 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c136
*+ bl_0_136 br_0_136 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c136
*+ bl_0_136 br_0_136 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c136
*+ bl_0_136 br_0_136 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c136
*+ bl_0_136 br_0_136 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c136
*+ bl_0_136 br_0_136 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c136
*+ bl_0_136 br_0_136 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c136
*+ bl_0_136 br_0_136 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c136
*+ bl_0_136 br_0_136 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c136
*+ bl_0_136 br_0_136 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c136
*+ bl_0_136 br_0_136 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c136
*+ bl_0_136 br_0_136 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c136
*+ bl_0_136 br_0_136 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c136
*+ bl_0_136 br_0_136 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c136
*+ bl_0_136 br_0_136 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c136
*+ bl_0_136 br_0_136 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c136
*+ bl_0_136 br_0_136 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c136
*+ bl_0_136 br_0_136 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c136
*+ bl_0_136 br_0_136 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c136
*+ bl_0_136 br_0_136 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c136
*+ bl_0_136 br_0_136 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c136
*+ bl_0_136 br_0_136 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c136
*+ bl_0_136 br_0_136 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c136
*+ bl_0_136 br_0_136 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c136
*+ bl_0_136 br_0_136 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c136
*+ bl_0_136 br_0_136 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c136
*+ bl_0_136 br_0_136 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c136
*+ bl_0_136 br_0_136 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c136
*+ bl_0_136 br_0_136 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c136
*+ bl_0_136 br_0_136 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c136
*+ bl_0_136 br_0_136 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c136
*+ bl_0_136 br_0_136 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c136
*+ bl_0_136 br_0_136 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c136
*+ bl_0_136 br_0_136 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c136
*+ bl_0_136 br_0_136 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c136
*+ bl_0_136 br_0_136 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c136
*+ bl_0_136 br_0_136 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c136
*+ bl_0_136 br_0_136 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c136
*+ bl_0_136 br_0_136 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c136
*+ bl_0_136 br_0_136 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c136
*+ bl_0_136 br_0_136 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c136
*+ bl_0_136 br_0_136 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c136
+ bl_0_136 br_0_136 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c137
+ bl_0_137 br_0_137 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c137
*+ bl_0_137 br_0_137 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c137
*+ bl_0_137 br_0_137 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c137
*+ bl_0_137 br_0_137 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c137
*+ bl_0_137 br_0_137 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c137
*+ bl_0_137 br_0_137 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c137
*+ bl_0_137 br_0_137 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c137
*+ bl_0_137 br_0_137 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c137
*+ bl_0_137 br_0_137 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c137
*+ bl_0_137 br_0_137 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c137
*+ bl_0_137 br_0_137 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c137
*+ bl_0_137 br_0_137 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c137
*+ bl_0_137 br_0_137 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c137
*+ bl_0_137 br_0_137 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c137
*+ bl_0_137 br_0_137 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c137
*+ bl_0_137 br_0_137 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c137
*+ bl_0_137 br_0_137 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c137
*+ bl_0_137 br_0_137 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c137
*+ bl_0_137 br_0_137 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c137
*+ bl_0_137 br_0_137 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c137
*+ bl_0_137 br_0_137 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c137
*+ bl_0_137 br_0_137 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c137
*+ bl_0_137 br_0_137 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c137
*+ bl_0_137 br_0_137 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c137
*+ bl_0_137 br_0_137 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c137
*+ bl_0_137 br_0_137 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c137
*+ bl_0_137 br_0_137 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c137
*+ bl_0_137 br_0_137 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c137
*+ bl_0_137 br_0_137 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c137
*+ bl_0_137 br_0_137 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c137
*+ bl_0_137 br_0_137 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c137
*+ bl_0_137 br_0_137 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c137
*+ bl_0_137 br_0_137 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c137
*+ bl_0_137 br_0_137 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c137
*+ bl_0_137 br_0_137 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c137
*+ bl_0_137 br_0_137 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c137
*+ bl_0_137 br_0_137 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c137
*+ bl_0_137 br_0_137 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c137
*+ bl_0_137 br_0_137 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c137
*+ bl_0_137 br_0_137 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c137
*+ bl_0_137 br_0_137 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c137
*+ bl_0_137 br_0_137 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c137
*+ bl_0_137 br_0_137 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c137
*+ bl_0_137 br_0_137 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c137
*+ bl_0_137 br_0_137 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c137
*+ bl_0_137 br_0_137 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c137
*+ bl_0_137 br_0_137 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c137
*+ bl_0_137 br_0_137 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c137
*+ bl_0_137 br_0_137 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c137
*+ bl_0_137 br_0_137 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c137
*+ bl_0_137 br_0_137 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c137
*+ bl_0_137 br_0_137 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c137
*+ bl_0_137 br_0_137 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c137
*+ bl_0_137 br_0_137 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c137
*+ bl_0_137 br_0_137 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c137
*+ bl_0_137 br_0_137 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c137
*+ bl_0_137 br_0_137 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c137
*+ bl_0_137 br_0_137 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c137
*+ bl_0_137 br_0_137 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c137
*+ bl_0_137 br_0_137 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c137
*+ bl_0_137 br_0_137 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c137
*+ bl_0_137 br_0_137 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c137
*+ bl_0_137 br_0_137 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c137
*+ bl_0_137 br_0_137 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c137
*+ bl_0_137 br_0_137 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c137
*+ bl_0_137 br_0_137 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c137
*+ bl_0_137 br_0_137 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c137
*+ bl_0_137 br_0_137 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c137
*+ bl_0_137 br_0_137 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c137
*+ bl_0_137 br_0_137 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c137
*+ bl_0_137 br_0_137 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c137
*+ bl_0_137 br_0_137 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c137
*+ bl_0_137 br_0_137 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c137
*+ bl_0_137 br_0_137 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c137
*+ bl_0_137 br_0_137 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c137
*+ bl_0_137 br_0_137 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c137
*+ bl_0_137 br_0_137 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c137
*+ bl_0_137 br_0_137 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c137
*+ bl_0_137 br_0_137 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c137
*+ bl_0_137 br_0_137 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c137
*+ bl_0_137 br_0_137 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c137
*+ bl_0_137 br_0_137 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c137
*+ bl_0_137 br_0_137 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c137
*+ bl_0_137 br_0_137 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c137
*+ bl_0_137 br_0_137 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c137
*+ bl_0_137 br_0_137 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c137
*+ bl_0_137 br_0_137 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c137
*+ bl_0_137 br_0_137 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c137
*+ bl_0_137 br_0_137 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c137
*+ bl_0_137 br_0_137 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c137
*+ bl_0_137 br_0_137 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c137
*+ bl_0_137 br_0_137 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c137
*+ bl_0_137 br_0_137 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c137
*+ bl_0_137 br_0_137 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c137
*+ bl_0_137 br_0_137 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c137
*+ bl_0_137 br_0_137 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c137
*+ bl_0_137 br_0_137 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c137
*+ bl_0_137 br_0_137 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c137
*+ bl_0_137 br_0_137 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c137
*+ bl_0_137 br_0_137 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c137
*+ bl_0_137 br_0_137 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c137
*+ bl_0_137 br_0_137 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c137
*+ bl_0_137 br_0_137 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c137
*+ bl_0_137 br_0_137 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c137
*+ bl_0_137 br_0_137 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c137
*+ bl_0_137 br_0_137 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c137
*+ bl_0_137 br_0_137 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c137
*+ bl_0_137 br_0_137 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c137
*+ bl_0_137 br_0_137 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c137
*+ bl_0_137 br_0_137 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c137
*+ bl_0_137 br_0_137 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c137
*+ bl_0_137 br_0_137 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c137
*+ bl_0_137 br_0_137 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c137
*+ bl_0_137 br_0_137 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c137
*+ bl_0_137 br_0_137 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c137
*+ bl_0_137 br_0_137 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c137
*+ bl_0_137 br_0_137 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c137
*+ bl_0_137 br_0_137 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c137
*+ bl_0_137 br_0_137 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c137
*+ bl_0_137 br_0_137 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c137
*+ bl_0_137 br_0_137 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c137
*+ bl_0_137 br_0_137 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c137
*+ bl_0_137 br_0_137 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c137
*+ bl_0_137 br_0_137 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c137
*+ bl_0_137 br_0_137 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c137
*+ bl_0_137 br_0_137 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c137
*+ bl_0_137 br_0_137 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c137
+ bl_0_137 br_0_137 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c138
+ bl_0_138 br_0_138 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c138
*+ bl_0_138 br_0_138 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c138
*+ bl_0_138 br_0_138 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c138
*+ bl_0_138 br_0_138 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c138
*+ bl_0_138 br_0_138 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c138
*+ bl_0_138 br_0_138 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c138
*+ bl_0_138 br_0_138 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c138
*+ bl_0_138 br_0_138 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c138
*+ bl_0_138 br_0_138 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c138
*+ bl_0_138 br_0_138 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c138
*+ bl_0_138 br_0_138 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c138
*+ bl_0_138 br_0_138 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c138
*+ bl_0_138 br_0_138 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c138
*+ bl_0_138 br_0_138 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c138
*+ bl_0_138 br_0_138 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c138
*+ bl_0_138 br_0_138 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c138
*+ bl_0_138 br_0_138 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c138
*+ bl_0_138 br_0_138 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c138
*+ bl_0_138 br_0_138 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c138
*+ bl_0_138 br_0_138 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c138
*+ bl_0_138 br_0_138 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c138
*+ bl_0_138 br_0_138 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c138
*+ bl_0_138 br_0_138 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c138
*+ bl_0_138 br_0_138 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c138
*+ bl_0_138 br_0_138 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c138
*+ bl_0_138 br_0_138 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c138
*+ bl_0_138 br_0_138 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c138
*+ bl_0_138 br_0_138 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c138
*+ bl_0_138 br_0_138 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c138
*+ bl_0_138 br_0_138 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c138
*+ bl_0_138 br_0_138 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c138
*+ bl_0_138 br_0_138 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c138
*+ bl_0_138 br_0_138 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c138
*+ bl_0_138 br_0_138 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c138
*+ bl_0_138 br_0_138 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c138
*+ bl_0_138 br_0_138 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c138
*+ bl_0_138 br_0_138 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c138
*+ bl_0_138 br_0_138 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c138
*+ bl_0_138 br_0_138 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c138
*+ bl_0_138 br_0_138 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c138
*+ bl_0_138 br_0_138 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c138
*+ bl_0_138 br_0_138 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c138
*+ bl_0_138 br_0_138 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c138
*+ bl_0_138 br_0_138 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c138
*+ bl_0_138 br_0_138 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c138
*+ bl_0_138 br_0_138 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c138
*+ bl_0_138 br_0_138 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c138
*+ bl_0_138 br_0_138 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c138
*+ bl_0_138 br_0_138 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c138
*+ bl_0_138 br_0_138 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c138
*+ bl_0_138 br_0_138 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c138
*+ bl_0_138 br_0_138 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c138
*+ bl_0_138 br_0_138 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c138
*+ bl_0_138 br_0_138 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c138
*+ bl_0_138 br_0_138 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c138
*+ bl_0_138 br_0_138 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c138
*+ bl_0_138 br_0_138 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c138
*+ bl_0_138 br_0_138 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c138
*+ bl_0_138 br_0_138 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c138
*+ bl_0_138 br_0_138 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c138
*+ bl_0_138 br_0_138 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c138
*+ bl_0_138 br_0_138 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c138
*+ bl_0_138 br_0_138 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c138
*+ bl_0_138 br_0_138 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c138
*+ bl_0_138 br_0_138 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c138
*+ bl_0_138 br_0_138 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c138
*+ bl_0_138 br_0_138 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c138
*+ bl_0_138 br_0_138 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c138
*+ bl_0_138 br_0_138 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c138
*+ bl_0_138 br_0_138 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c138
*+ bl_0_138 br_0_138 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c138
*+ bl_0_138 br_0_138 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c138
*+ bl_0_138 br_0_138 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c138
*+ bl_0_138 br_0_138 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c138
*+ bl_0_138 br_0_138 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c138
*+ bl_0_138 br_0_138 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c138
*+ bl_0_138 br_0_138 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c138
*+ bl_0_138 br_0_138 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c138
*+ bl_0_138 br_0_138 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c138
*+ bl_0_138 br_0_138 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c138
*+ bl_0_138 br_0_138 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c138
*+ bl_0_138 br_0_138 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c138
*+ bl_0_138 br_0_138 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c138
*+ bl_0_138 br_0_138 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c138
*+ bl_0_138 br_0_138 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c138
*+ bl_0_138 br_0_138 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c138
*+ bl_0_138 br_0_138 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c138
*+ bl_0_138 br_0_138 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c138
*+ bl_0_138 br_0_138 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c138
*+ bl_0_138 br_0_138 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c138
*+ bl_0_138 br_0_138 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c138
*+ bl_0_138 br_0_138 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c138
*+ bl_0_138 br_0_138 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c138
*+ bl_0_138 br_0_138 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c138
*+ bl_0_138 br_0_138 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c138
*+ bl_0_138 br_0_138 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c138
*+ bl_0_138 br_0_138 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c138
*+ bl_0_138 br_0_138 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c138
*+ bl_0_138 br_0_138 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c138
*+ bl_0_138 br_0_138 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c138
*+ bl_0_138 br_0_138 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c138
*+ bl_0_138 br_0_138 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c138
*+ bl_0_138 br_0_138 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c138
*+ bl_0_138 br_0_138 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c138
*+ bl_0_138 br_0_138 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c138
*+ bl_0_138 br_0_138 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c138
*+ bl_0_138 br_0_138 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c138
*+ bl_0_138 br_0_138 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c138
*+ bl_0_138 br_0_138 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c138
*+ bl_0_138 br_0_138 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c138
*+ bl_0_138 br_0_138 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c138
*+ bl_0_138 br_0_138 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c138
*+ bl_0_138 br_0_138 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c138
*+ bl_0_138 br_0_138 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c138
*+ bl_0_138 br_0_138 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c138
*+ bl_0_138 br_0_138 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c138
*+ bl_0_138 br_0_138 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c138
*+ bl_0_138 br_0_138 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c138
*+ bl_0_138 br_0_138 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c138
*+ bl_0_138 br_0_138 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c138
*+ bl_0_138 br_0_138 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c138
*+ bl_0_138 br_0_138 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c138
*+ bl_0_138 br_0_138 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c138
*+ bl_0_138 br_0_138 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c138
*+ bl_0_138 br_0_138 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c138
*+ bl_0_138 br_0_138 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c138
*+ bl_0_138 br_0_138 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c138
+ bl_0_138 br_0_138 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c139
+ bl_0_139 br_0_139 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c139
*+ bl_0_139 br_0_139 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c139
*+ bl_0_139 br_0_139 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c139
*+ bl_0_139 br_0_139 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c139
*+ bl_0_139 br_0_139 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c139
*+ bl_0_139 br_0_139 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c139
*+ bl_0_139 br_0_139 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c139
*+ bl_0_139 br_0_139 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c139
*+ bl_0_139 br_0_139 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c139
*+ bl_0_139 br_0_139 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c139
*+ bl_0_139 br_0_139 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c139
*+ bl_0_139 br_0_139 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c139
*+ bl_0_139 br_0_139 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c139
*+ bl_0_139 br_0_139 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c139
*+ bl_0_139 br_0_139 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c139
*+ bl_0_139 br_0_139 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c139
*+ bl_0_139 br_0_139 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c139
*+ bl_0_139 br_0_139 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c139
*+ bl_0_139 br_0_139 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c139
*+ bl_0_139 br_0_139 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c139
*+ bl_0_139 br_0_139 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c139
*+ bl_0_139 br_0_139 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c139
*+ bl_0_139 br_0_139 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c139
*+ bl_0_139 br_0_139 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c139
*+ bl_0_139 br_0_139 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c139
*+ bl_0_139 br_0_139 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c139
*+ bl_0_139 br_0_139 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c139
*+ bl_0_139 br_0_139 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c139
*+ bl_0_139 br_0_139 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c139
*+ bl_0_139 br_0_139 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c139
*+ bl_0_139 br_0_139 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c139
*+ bl_0_139 br_0_139 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c139
*+ bl_0_139 br_0_139 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c139
*+ bl_0_139 br_0_139 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c139
*+ bl_0_139 br_0_139 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c139
*+ bl_0_139 br_0_139 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c139
*+ bl_0_139 br_0_139 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c139
*+ bl_0_139 br_0_139 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c139
*+ bl_0_139 br_0_139 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c139
*+ bl_0_139 br_0_139 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c139
*+ bl_0_139 br_0_139 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c139
*+ bl_0_139 br_0_139 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c139
*+ bl_0_139 br_0_139 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c139
*+ bl_0_139 br_0_139 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c139
*+ bl_0_139 br_0_139 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c139
*+ bl_0_139 br_0_139 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c139
*+ bl_0_139 br_0_139 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c139
*+ bl_0_139 br_0_139 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c139
*+ bl_0_139 br_0_139 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c139
*+ bl_0_139 br_0_139 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c139
*+ bl_0_139 br_0_139 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c139
*+ bl_0_139 br_0_139 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c139
*+ bl_0_139 br_0_139 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c139
*+ bl_0_139 br_0_139 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c139
*+ bl_0_139 br_0_139 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c139
*+ bl_0_139 br_0_139 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c139
*+ bl_0_139 br_0_139 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c139
*+ bl_0_139 br_0_139 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c139
*+ bl_0_139 br_0_139 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c139
*+ bl_0_139 br_0_139 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c139
*+ bl_0_139 br_0_139 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c139
*+ bl_0_139 br_0_139 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c139
*+ bl_0_139 br_0_139 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c139
*+ bl_0_139 br_0_139 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c139
*+ bl_0_139 br_0_139 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c139
*+ bl_0_139 br_0_139 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c139
*+ bl_0_139 br_0_139 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c139
*+ bl_0_139 br_0_139 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c139
*+ bl_0_139 br_0_139 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c139
*+ bl_0_139 br_0_139 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c139
*+ bl_0_139 br_0_139 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c139
*+ bl_0_139 br_0_139 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c139
*+ bl_0_139 br_0_139 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c139
*+ bl_0_139 br_0_139 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c139
*+ bl_0_139 br_0_139 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c139
*+ bl_0_139 br_0_139 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c139
*+ bl_0_139 br_0_139 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c139
*+ bl_0_139 br_0_139 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c139
*+ bl_0_139 br_0_139 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c139
*+ bl_0_139 br_0_139 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c139
*+ bl_0_139 br_0_139 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c139
*+ bl_0_139 br_0_139 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c139
*+ bl_0_139 br_0_139 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c139
*+ bl_0_139 br_0_139 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c139
*+ bl_0_139 br_0_139 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c139
*+ bl_0_139 br_0_139 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c139
*+ bl_0_139 br_0_139 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c139
*+ bl_0_139 br_0_139 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c139
*+ bl_0_139 br_0_139 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c139
*+ bl_0_139 br_0_139 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c139
*+ bl_0_139 br_0_139 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c139
*+ bl_0_139 br_0_139 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c139
*+ bl_0_139 br_0_139 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c139
*+ bl_0_139 br_0_139 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c139
*+ bl_0_139 br_0_139 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c139
*+ bl_0_139 br_0_139 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c139
*+ bl_0_139 br_0_139 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c139
*+ bl_0_139 br_0_139 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c139
*+ bl_0_139 br_0_139 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c139
*+ bl_0_139 br_0_139 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c139
*+ bl_0_139 br_0_139 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c139
*+ bl_0_139 br_0_139 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c139
*+ bl_0_139 br_0_139 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c139
*+ bl_0_139 br_0_139 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c139
*+ bl_0_139 br_0_139 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c139
*+ bl_0_139 br_0_139 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c139
*+ bl_0_139 br_0_139 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c139
*+ bl_0_139 br_0_139 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c139
*+ bl_0_139 br_0_139 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c139
*+ bl_0_139 br_0_139 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c139
*+ bl_0_139 br_0_139 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c139
*+ bl_0_139 br_0_139 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c139
*+ bl_0_139 br_0_139 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c139
*+ bl_0_139 br_0_139 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c139
*+ bl_0_139 br_0_139 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c139
*+ bl_0_139 br_0_139 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c139
*+ bl_0_139 br_0_139 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c139
*+ bl_0_139 br_0_139 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c139
*+ bl_0_139 br_0_139 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c139
*+ bl_0_139 br_0_139 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c139
*+ bl_0_139 br_0_139 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c139
*+ bl_0_139 br_0_139 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c139
*+ bl_0_139 br_0_139 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c139
*+ bl_0_139 br_0_139 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c139
*+ bl_0_139 br_0_139 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c139
*+ bl_0_139 br_0_139 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c139
*+ bl_0_139 br_0_139 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c139
+ bl_0_139 br_0_139 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c140
+ bl_0_140 br_0_140 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c140
*+ bl_0_140 br_0_140 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c140
*+ bl_0_140 br_0_140 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c140
*+ bl_0_140 br_0_140 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c140
*+ bl_0_140 br_0_140 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c140
*+ bl_0_140 br_0_140 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c140
*+ bl_0_140 br_0_140 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c140
*+ bl_0_140 br_0_140 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c140
*+ bl_0_140 br_0_140 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c140
*+ bl_0_140 br_0_140 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c140
*+ bl_0_140 br_0_140 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c140
*+ bl_0_140 br_0_140 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c140
*+ bl_0_140 br_0_140 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c140
*+ bl_0_140 br_0_140 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c140
*+ bl_0_140 br_0_140 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c140
*+ bl_0_140 br_0_140 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c140
*+ bl_0_140 br_0_140 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c140
*+ bl_0_140 br_0_140 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c140
*+ bl_0_140 br_0_140 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c140
*+ bl_0_140 br_0_140 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c140
*+ bl_0_140 br_0_140 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c140
*+ bl_0_140 br_0_140 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c140
*+ bl_0_140 br_0_140 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c140
*+ bl_0_140 br_0_140 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c140
*+ bl_0_140 br_0_140 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c140
*+ bl_0_140 br_0_140 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c140
*+ bl_0_140 br_0_140 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c140
*+ bl_0_140 br_0_140 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c140
*+ bl_0_140 br_0_140 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c140
*+ bl_0_140 br_0_140 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c140
*+ bl_0_140 br_0_140 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c140
*+ bl_0_140 br_0_140 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c140
*+ bl_0_140 br_0_140 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c140
*+ bl_0_140 br_0_140 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c140
*+ bl_0_140 br_0_140 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c140
*+ bl_0_140 br_0_140 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c140
*+ bl_0_140 br_0_140 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c140
*+ bl_0_140 br_0_140 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c140
*+ bl_0_140 br_0_140 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c140
*+ bl_0_140 br_0_140 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c140
*+ bl_0_140 br_0_140 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c140
*+ bl_0_140 br_0_140 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c140
*+ bl_0_140 br_0_140 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c140
*+ bl_0_140 br_0_140 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c140
*+ bl_0_140 br_0_140 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c140
*+ bl_0_140 br_0_140 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c140
*+ bl_0_140 br_0_140 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c140
*+ bl_0_140 br_0_140 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c140
*+ bl_0_140 br_0_140 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c140
*+ bl_0_140 br_0_140 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c140
*+ bl_0_140 br_0_140 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c140
*+ bl_0_140 br_0_140 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c140
*+ bl_0_140 br_0_140 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c140
*+ bl_0_140 br_0_140 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c140
*+ bl_0_140 br_0_140 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c140
*+ bl_0_140 br_0_140 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c140
*+ bl_0_140 br_0_140 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c140
*+ bl_0_140 br_0_140 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c140
*+ bl_0_140 br_0_140 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c140
*+ bl_0_140 br_0_140 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c140
*+ bl_0_140 br_0_140 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c140
*+ bl_0_140 br_0_140 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c140
*+ bl_0_140 br_0_140 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c140
*+ bl_0_140 br_0_140 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c140
*+ bl_0_140 br_0_140 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c140
*+ bl_0_140 br_0_140 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c140
*+ bl_0_140 br_0_140 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c140
*+ bl_0_140 br_0_140 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c140
*+ bl_0_140 br_0_140 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c140
*+ bl_0_140 br_0_140 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c140
*+ bl_0_140 br_0_140 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c140
*+ bl_0_140 br_0_140 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c140
*+ bl_0_140 br_0_140 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c140
*+ bl_0_140 br_0_140 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c140
*+ bl_0_140 br_0_140 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c140
*+ bl_0_140 br_0_140 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c140
*+ bl_0_140 br_0_140 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c140
*+ bl_0_140 br_0_140 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c140
*+ bl_0_140 br_0_140 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c140
*+ bl_0_140 br_0_140 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c140
*+ bl_0_140 br_0_140 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c140
*+ bl_0_140 br_0_140 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c140
*+ bl_0_140 br_0_140 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c140
*+ bl_0_140 br_0_140 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c140
*+ bl_0_140 br_0_140 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c140
*+ bl_0_140 br_0_140 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c140
*+ bl_0_140 br_0_140 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c140
*+ bl_0_140 br_0_140 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c140
*+ bl_0_140 br_0_140 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c140
*+ bl_0_140 br_0_140 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c140
*+ bl_0_140 br_0_140 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c140
*+ bl_0_140 br_0_140 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c140
*+ bl_0_140 br_0_140 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c140
*+ bl_0_140 br_0_140 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c140
*+ bl_0_140 br_0_140 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c140
*+ bl_0_140 br_0_140 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c140
*+ bl_0_140 br_0_140 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c140
*+ bl_0_140 br_0_140 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c140
*+ bl_0_140 br_0_140 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c140
*+ bl_0_140 br_0_140 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c140
*+ bl_0_140 br_0_140 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c140
*+ bl_0_140 br_0_140 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c140
*+ bl_0_140 br_0_140 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c140
*+ bl_0_140 br_0_140 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c140
*+ bl_0_140 br_0_140 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c140
*+ bl_0_140 br_0_140 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c140
*+ bl_0_140 br_0_140 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c140
*+ bl_0_140 br_0_140 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c140
*+ bl_0_140 br_0_140 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c140
*+ bl_0_140 br_0_140 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c140
*+ bl_0_140 br_0_140 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c140
*+ bl_0_140 br_0_140 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c140
*+ bl_0_140 br_0_140 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c140
*+ bl_0_140 br_0_140 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c140
*+ bl_0_140 br_0_140 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c140
*+ bl_0_140 br_0_140 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c140
*+ bl_0_140 br_0_140 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c140
*+ bl_0_140 br_0_140 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c140
*+ bl_0_140 br_0_140 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c140
*+ bl_0_140 br_0_140 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c140
*+ bl_0_140 br_0_140 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c140
*+ bl_0_140 br_0_140 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c140
*+ bl_0_140 br_0_140 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c140
*+ bl_0_140 br_0_140 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c140
*+ bl_0_140 br_0_140 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c140
*+ bl_0_140 br_0_140 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c140
*+ bl_0_140 br_0_140 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c140
+ bl_0_140 br_0_140 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c141
+ bl_0_141 br_0_141 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c141
*+ bl_0_141 br_0_141 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c141
*+ bl_0_141 br_0_141 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c141
*+ bl_0_141 br_0_141 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c141
*+ bl_0_141 br_0_141 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c141
*+ bl_0_141 br_0_141 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c141
*+ bl_0_141 br_0_141 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c141
*+ bl_0_141 br_0_141 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c141
*+ bl_0_141 br_0_141 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c141
*+ bl_0_141 br_0_141 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c141
*+ bl_0_141 br_0_141 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c141
*+ bl_0_141 br_0_141 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c141
*+ bl_0_141 br_0_141 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c141
*+ bl_0_141 br_0_141 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c141
*+ bl_0_141 br_0_141 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c141
*+ bl_0_141 br_0_141 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c141
*+ bl_0_141 br_0_141 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c141
*+ bl_0_141 br_0_141 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c141
*+ bl_0_141 br_0_141 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c141
*+ bl_0_141 br_0_141 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c141
*+ bl_0_141 br_0_141 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c141
*+ bl_0_141 br_0_141 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c141
*+ bl_0_141 br_0_141 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c141
*+ bl_0_141 br_0_141 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c141
*+ bl_0_141 br_0_141 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c141
*+ bl_0_141 br_0_141 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c141
*+ bl_0_141 br_0_141 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c141
*+ bl_0_141 br_0_141 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c141
*+ bl_0_141 br_0_141 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c141
*+ bl_0_141 br_0_141 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c141
*+ bl_0_141 br_0_141 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c141
*+ bl_0_141 br_0_141 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c141
*+ bl_0_141 br_0_141 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c141
*+ bl_0_141 br_0_141 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c141
*+ bl_0_141 br_0_141 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c141
*+ bl_0_141 br_0_141 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c141
*+ bl_0_141 br_0_141 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c141
*+ bl_0_141 br_0_141 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c141
*+ bl_0_141 br_0_141 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c141
*+ bl_0_141 br_0_141 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c141
*+ bl_0_141 br_0_141 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c141
*+ bl_0_141 br_0_141 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c141
*+ bl_0_141 br_0_141 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c141
*+ bl_0_141 br_0_141 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c141
*+ bl_0_141 br_0_141 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c141
*+ bl_0_141 br_0_141 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c141
*+ bl_0_141 br_0_141 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c141
*+ bl_0_141 br_0_141 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c141
*+ bl_0_141 br_0_141 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c141
*+ bl_0_141 br_0_141 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c141
*+ bl_0_141 br_0_141 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c141
*+ bl_0_141 br_0_141 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c141
*+ bl_0_141 br_0_141 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c141
*+ bl_0_141 br_0_141 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c141
*+ bl_0_141 br_0_141 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c141
*+ bl_0_141 br_0_141 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c141
*+ bl_0_141 br_0_141 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c141
*+ bl_0_141 br_0_141 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c141
*+ bl_0_141 br_0_141 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c141
*+ bl_0_141 br_0_141 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c141
*+ bl_0_141 br_0_141 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c141
*+ bl_0_141 br_0_141 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c141
*+ bl_0_141 br_0_141 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c141
*+ bl_0_141 br_0_141 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c141
*+ bl_0_141 br_0_141 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c141
*+ bl_0_141 br_0_141 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c141
*+ bl_0_141 br_0_141 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c141
*+ bl_0_141 br_0_141 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c141
*+ bl_0_141 br_0_141 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c141
*+ bl_0_141 br_0_141 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c141
*+ bl_0_141 br_0_141 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c141
*+ bl_0_141 br_0_141 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c141
*+ bl_0_141 br_0_141 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c141
*+ bl_0_141 br_0_141 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c141
*+ bl_0_141 br_0_141 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c141
*+ bl_0_141 br_0_141 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c141
*+ bl_0_141 br_0_141 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c141
*+ bl_0_141 br_0_141 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c141
*+ bl_0_141 br_0_141 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c141
*+ bl_0_141 br_0_141 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c141
*+ bl_0_141 br_0_141 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c141
*+ bl_0_141 br_0_141 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c141
*+ bl_0_141 br_0_141 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c141
*+ bl_0_141 br_0_141 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c141
*+ bl_0_141 br_0_141 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c141
*+ bl_0_141 br_0_141 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c141
*+ bl_0_141 br_0_141 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c141
*+ bl_0_141 br_0_141 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c141
*+ bl_0_141 br_0_141 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c141
*+ bl_0_141 br_0_141 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c141
*+ bl_0_141 br_0_141 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c141
*+ bl_0_141 br_0_141 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c141
*+ bl_0_141 br_0_141 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c141
*+ bl_0_141 br_0_141 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c141
*+ bl_0_141 br_0_141 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c141
*+ bl_0_141 br_0_141 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c141
*+ bl_0_141 br_0_141 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c141
*+ bl_0_141 br_0_141 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c141
*+ bl_0_141 br_0_141 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c141
*+ bl_0_141 br_0_141 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c141
*+ bl_0_141 br_0_141 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c141
*+ bl_0_141 br_0_141 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c141
*+ bl_0_141 br_0_141 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c141
*+ bl_0_141 br_0_141 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c141
*+ bl_0_141 br_0_141 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c141
*+ bl_0_141 br_0_141 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c141
*+ bl_0_141 br_0_141 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c141
*+ bl_0_141 br_0_141 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c141
*+ bl_0_141 br_0_141 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c141
*+ bl_0_141 br_0_141 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c141
*+ bl_0_141 br_0_141 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c141
*+ bl_0_141 br_0_141 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c141
*+ bl_0_141 br_0_141 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c141
*+ bl_0_141 br_0_141 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c141
*+ bl_0_141 br_0_141 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c141
*+ bl_0_141 br_0_141 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c141
*+ bl_0_141 br_0_141 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c141
*+ bl_0_141 br_0_141 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c141
*+ bl_0_141 br_0_141 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c141
*+ bl_0_141 br_0_141 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c141
*+ bl_0_141 br_0_141 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c141
*+ bl_0_141 br_0_141 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c141
*+ bl_0_141 br_0_141 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c141
*+ bl_0_141 br_0_141 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c141
*+ bl_0_141 br_0_141 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c141
*+ bl_0_141 br_0_141 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c141
*+ bl_0_141 br_0_141 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c141
+ bl_0_141 br_0_141 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c142
+ bl_0_142 br_0_142 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c142
*+ bl_0_142 br_0_142 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c142
*+ bl_0_142 br_0_142 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c142
*+ bl_0_142 br_0_142 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c142
*+ bl_0_142 br_0_142 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c142
*+ bl_0_142 br_0_142 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c142
*+ bl_0_142 br_0_142 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c142
*+ bl_0_142 br_0_142 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c142
*+ bl_0_142 br_0_142 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c142
*+ bl_0_142 br_0_142 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c142
*+ bl_0_142 br_0_142 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c142
*+ bl_0_142 br_0_142 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c142
*+ bl_0_142 br_0_142 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c142
*+ bl_0_142 br_0_142 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c142
*+ bl_0_142 br_0_142 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c142
*+ bl_0_142 br_0_142 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c142
*+ bl_0_142 br_0_142 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c142
*+ bl_0_142 br_0_142 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c142
*+ bl_0_142 br_0_142 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c142
*+ bl_0_142 br_0_142 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c142
*+ bl_0_142 br_0_142 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c142
*+ bl_0_142 br_0_142 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c142
*+ bl_0_142 br_0_142 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c142
*+ bl_0_142 br_0_142 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c142
*+ bl_0_142 br_0_142 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c142
*+ bl_0_142 br_0_142 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c142
*+ bl_0_142 br_0_142 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c142
*+ bl_0_142 br_0_142 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c142
*+ bl_0_142 br_0_142 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c142
*+ bl_0_142 br_0_142 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c142
*+ bl_0_142 br_0_142 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c142
*+ bl_0_142 br_0_142 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c142
*+ bl_0_142 br_0_142 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c142
*+ bl_0_142 br_0_142 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c142
*+ bl_0_142 br_0_142 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c142
*+ bl_0_142 br_0_142 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c142
*+ bl_0_142 br_0_142 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c142
*+ bl_0_142 br_0_142 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c142
*+ bl_0_142 br_0_142 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c142
*+ bl_0_142 br_0_142 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c142
*+ bl_0_142 br_0_142 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c142
*+ bl_0_142 br_0_142 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c142
*+ bl_0_142 br_0_142 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c142
*+ bl_0_142 br_0_142 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c142
*+ bl_0_142 br_0_142 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c142
*+ bl_0_142 br_0_142 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c142
*+ bl_0_142 br_0_142 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c142
*+ bl_0_142 br_0_142 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c142
*+ bl_0_142 br_0_142 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c142
*+ bl_0_142 br_0_142 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c142
*+ bl_0_142 br_0_142 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c142
*+ bl_0_142 br_0_142 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c142
*+ bl_0_142 br_0_142 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c142
*+ bl_0_142 br_0_142 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c142
*+ bl_0_142 br_0_142 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c142
*+ bl_0_142 br_0_142 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c142
*+ bl_0_142 br_0_142 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c142
*+ bl_0_142 br_0_142 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c142
*+ bl_0_142 br_0_142 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c142
*+ bl_0_142 br_0_142 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c142
*+ bl_0_142 br_0_142 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c142
*+ bl_0_142 br_0_142 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c142
*+ bl_0_142 br_0_142 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c142
*+ bl_0_142 br_0_142 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c142
*+ bl_0_142 br_0_142 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c142
*+ bl_0_142 br_0_142 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c142
*+ bl_0_142 br_0_142 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c142
*+ bl_0_142 br_0_142 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c142
*+ bl_0_142 br_0_142 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c142
*+ bl_0_142 br_0_142 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c142
*+ bl_0_142 br_0_142 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c142
*+ bl_0_142 br_0_142 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c142
*+ bl_0_142 br_0_142 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c142
*+ bl_0_142 br_0_142 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c142
*+ bl_0_142 br_0_142 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c142
*+ bl_0_142 br_0_142 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c142
*+ bl_0_142 br_0_142 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c142
*+ bl_0_142 br_0_142 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c142
*+ bl_0_142 br_0_142 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c142
*+ bl_0_142 br_0_142 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c142
*+ bl_0_142 br_0_142 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c142
*+ bl_0_142 br_0_142 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c142
*+ bl_0_142 br_0_142 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c142
*+ bl_0_142 br_0_142 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c142
*+ bl_0_142 br_0_142 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c142
*+ bl_0_142 br_0_142 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c142
*+ bl_0_142 br_0_142 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c142
*+ bl_0_142 br_0_142 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c142
*+ bl_0_142 br_0_142 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c142
*+ bl_0_142 br_0_142 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c142
*+ bl_0_142 br_0_142 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c142
*+ bl_0_142 br_0_142 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c142
*+ bl_0_142 br_0_142 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c142
*+ bl_0_142 br_0_142 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c142
*+ bl_0_142 br_0_142 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c142
*+ bl_0_142 br_0_142 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c142
*+ bl_0_142 br_0_142 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c142
*+ bl_0_142 br_0_142 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c142
*+ bl_0_142 br_0_142 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c142
*+ bl_0_142 br_0_142 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c142
*+ bl_0_142 br_0_142 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c142
*+ bl_0_142 br_0_142 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c142
*+ bl_0_142 br_0_142 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c142
*+ bl_0_142 br_0_142 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c142
*+ bl_0_142 br_0_142 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c142
*+ bl_0_142 br_0_142 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c142
*+ bl_0_142 br_0_142 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c142
*+ bl_0_142 br_0_142 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c142
*+ bl_0_142 br_0_142 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c142
*+ bl_0_142 br_0_142 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c142
*+ bl_0_142 br_0_142 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c142
*+ bl_0_142 br_0_142 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c142
*+ bl_0_142 br_0_142 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c142
*+ bl_0_142 br_0_142 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c142
*+ bl_0_142 br_0_142 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c142
*+ bl_0_142 br_0_142 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c142
*+ bl_0_142 br_0_142 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c142
*+ bl_0_142 br_0_142 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c142
*+ bl_0_142 br_0_142 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c142
*+ bl_0_142 br_0_142 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c142
*+ bl_0_142 br_0_142 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c142
*+ bl_0_142 br_0_142 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c142
*+ bl_0_142 br_0_142 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c142
*+ bl_0_142 br_0_142 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c142
*+ bl_0_142 br_0_142 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c142
*+ bl_0_142 br_0_142 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c142
*+ bl_0_142 br_0_142 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c142
+ bl_0_142 br_0_142 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c143
+ bl_0_143 br_0_143 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c143
*+ bl_0_143 br_0_143 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c143
*+ bl_0_143 br_0_143 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c143
*+ bl_0_143 br_0_143 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c143
*+ bl_0_143 br_0_143 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c143
*+ bl_0_143 br_0_143 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c143
*+ bl_0_143 br_0_143 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c143
*+ bl_0_143 br_0_143 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c143
*+ bl_0_143 br_0_143 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c143
*+ bl_0_143 br_0_143 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c143
*+ bl_0_143 br_0_143 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c143
*+ bl_0_143 br_0_143 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c143
*+ bl_0_143 br_0_143 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c143
*+ bl_0_143 br_0_143 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c143
*+ bl_0_143 br_0_143 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c143
*+ bl_0_143 br_0_143 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c143
*+ bl_0_143 br_0_143 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c143
*+ bl_0_143 br_0_143 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c143
*+ bl_0_143 br_0_143 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c143
*+ bl_0_143 br_0_143 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c143
*+ bl_0_143 br_0_143 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c143
*+ bl_0_143 br_0_143 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c143
*+ bl_0_143 br_0_143 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c143
*+ bl_0_143 br_0_143 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c143
*+ bl_0_143 br_0_143 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c143
*+ bl_0_143 br_0_143 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c143
*+ bl_0_143 br_0_143 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c143
*+ bl_0_143 br_0_143 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c143
*+ bl_0_143 br_0_143 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c143
*+ bl_0_143 br_0_143 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c143
*+ bl_0_143 br_0_143 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c143
*+ bl_0_143 br_0_143 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c143
*+ bl_0_143 br_0_143 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c143
*+ bl_0_143 br_0_143 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c143
*+ bl_0_143 br_0_143 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c143
*+ bl_0_143 br_0_143 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c143
*+ bl_0_143 br_0_143 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c143
*+ bl_0_143 br_0_143 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c143
*+ bl_0_143 br_0_143 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c143
*+ bl_0_143 br_0_143 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c143
*+ bl_0_143 br_0_143 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c143
*+ bl_0_143 br_0_143 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c143
*+ bl_0_143 br_0_143 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c143
*+ bl_0_143 br_0_143 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c143
*+ bl_0_143 br_0_143 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c143
*+ bl_0_143 br_0_143 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c143
*+ bl_0_143 br_0_143 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c143
*+ bl_0_143 br_0_143 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c143
*+ bl_0_143 br_0_143 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c143
*+ bl_0_143 br_0_143 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c143
*+ bl_0_143 br_0_143 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c143
*+ bl_0_143 br_0_143 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c143
*+ bl_0_143 br_0_143 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c143
*+ bl_0_143 br_0_143 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c143
*+ bl_0_143 br_0_143 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c143
*+ bl_0_143 br_0_143 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c143
*+ bl_0_143 br_0_143 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c143
*+ bl_0_143 br_0_143 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c143
*+ bl_0_143 br_0_143 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c143
*+ bl_0_143 br_0_143 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c143
*+ bl_0_143 br_0_143 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c143
*+ bl_0_143 br_0_143 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c143
*+ bl_0_143 br_0_143 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c143
*+ bl_0_143 br_0_143 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c143
*+ bl_0_143 br_0_143 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c143
*+ bl_0_143 br_0_143 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c143
*+ bl_0_143 br_0_143 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c143
*+ bl_0_143 br_0_143 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c143
*+ bl_0_143 br_0_143 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c143
*+ bl_0_143 br_0_143 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c143
*+ bl_0_143 br_0_143 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c143
*+ bl_0_143 br_0_143 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c143
*+ bl_0_143 br_0_143 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c143
*+ bl_0_143 br_0_143 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c143
*+ bl_0_143 br_0_143 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c143
*+ bl_0_143 br_0_143 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c143
*+ bl_0_143 br_0_143 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c143
*+ bl_0_143 br_0_143 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c143
*+ bl_0_143 br_0_143 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c143
*+ bl_0_143 br_0_143 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c143
*+ bl_0_143 br_0_143 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c143
*+ bl_0_143 br_0_143 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c143
*+ bl_0_143 br_0_143 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c143
*+ bl_0_143 br_0_143 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c143
*+ bl_0_143 br_0_143 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c143
*+ bl_0_143 br_0_143 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c143
*+ bl_0_143 br_0_143 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c143
*+ bl_0_143 br_0_143 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c143
*+ bl_0_143 br_0_143 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c143
*+ bl_0_143 br_0_143 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c143
*+ bl_0_143 br_0_143 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c143
*+ bl_0_143 br_0_143 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c143
*+ bl_0_143 br_0_143 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c143
*+ bl_0_143 br_0_143 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c143
*+ bl_0_143 br_0_143 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c143
*+ bl_0_143 br_0_143 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c143
*+ bl_0_143 br_0_143 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c143
*+ bl_0_143 br_0_143 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c143
*+ bl_0_143 br_0_143 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c143
*+ bl_0_143 br_0_143 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c143
*+ bl_0_143 br_0_143 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c143
*+ bl_0_143 br_0_143 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c143
*+ bl_0_143 br_0_143 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c143
*+ bl_0_143 br_0_143 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c143
*+ bl_0_143 br_0_143 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c143
*+ bl_0_143 br_0_143 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c143
*+ bl_0_143 br_0_143 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c143
*+ bl_0_143 br_0_143 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c143
*+ bl_0_143 br_0_143 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c143
*+ bl_0_143 br_0_143 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c143
*+ bl_0_143 br_0_143 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c143
*+ bl_0_143 br_0_143 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c143
*+ bl_0_143 br_0_143 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c143
*+ bl_0_143 br_0_143 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c143
*+ bl_0_143 br_0_143 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c143
*+ bl_0_143 br_0_143 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c143
*+ bl_0_143 br_0_143 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c143
*+ bl_0_143 br_0_143 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c143
*+ bl_0_143 br_0_143 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c143
*+ bl_0_143 br_0_143 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c143
*+ bl_0_143 br_0_143 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c143
*+ bl_0_143 br_0_143 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c143
*+ bl_0_143 br_0_143 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c143
*+ bl_0_143 br_0_143 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c143
*+ bl_0_143 br_0_143 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c143
*+ bl_0_143 br_0_143 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c143
*+ bl_0_143 br_0_143 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c143
+ bl_0_143 br_0_143 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c144
+ bl_0_144 br_0_144 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c144
*+ bl_0_144 br_0_144 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c144
*+ bl_0_144 br_0_144 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c144
*+ bl_0_144 br_0_144 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c144
*+ bl_0_144 br_0_144 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c144
*+ bl_0_144 br_0_144 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c144
*+ bl_0_144 br_0_144 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c144
*+ bl_0_144 br_0_144 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c144
*+ bl_0_144 br_0_144 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c144
*+ bl_0_144 br_0_144 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c144
*+ bl_0_144 br_0_144 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c144
*+ bl_0_144 br_0_144 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c144
*+ bl_0_144 br_0_144 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c144
*+ bl_0_144 br_0_144 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c144
*+ bl_0_144 br_0_144 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c144
*+ bl_0_144 br_0_144 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c144
*+ bl_0_144 br_0_144 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c144
*+ bl_0_144 br_0_144 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c144
*+ bl_0_144 br_0_144 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c144
*+ bl_0_144 br_0_144 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c144
*+ bl_0_144 br_0_144 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c144
*+ bl_0_144 br_0_144 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c144
*+ bl_0_144 br_0_144 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c144
*+ bl_0_144 br_0_144 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c144
*+ bl_0_144 br_0_144 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c144
*+ bl_0_144 br_0_144 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c144
*+ bl_0_144 br_0_144 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c144
*+ bl_0_144 br_0_144 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c144
*+ bl_0_144 br_0_144 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c144
*+ bl_0_144 br_0_144 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c144
*+ bl_0_144 br_0_144 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c144
*+ bl_0_144 br_0_144 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c144
*+ bl_0_144 br_0_144 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c144
*+ bl_0_144 br_0_144 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c144
*+ bl_0_144 br_0_144 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c144
*+ bl_0_144 br_0_144 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c144
*+ bl_0_144 br_0_144 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c144
*+ bl_0_144 br_0_144 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c144
*+ bl_0_144 br_0_144 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c144
*+ bl_0_144 br_0_144 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c144
*+ bl_0_144 br_0_144 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c144
*+ bl_0_144 br_0_144 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c144
*+ bl_0_144 br_0_144 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c144
*+ bl_0_144 br_0_144 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c144
*+ bl_0_144 br_0_144 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c144
*+ bl_0_144 br_0_144 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c144
*+ bl_0_144 br_0_144 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c144
*+ bl_0_144 br_0_144 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c144
*+ bl_0_144 br_0_144 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c144
*+ bl_0_144 br_0_144 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c144
*+ bl_0_144 br_0_144 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c144
*+ bl_0_144 br_0_144 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c144
*+ bl_0_144 br_0_144 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c144
*+ bl_0_144 br_0_144 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c144
*+ bl_0_144 br_0_144 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c144
*+ bl_0_144 br_0_144 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c144
*+ bl_0_144 br_0_144 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c144
*+ bl_0_144 br_0_144 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c144
*+ bl_0_144 br_0_144 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c144
*+ bl_0_144 br_0_144 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c144
*+ bl_0_144 br_0_144 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c144
*+ bl_0_144 br_0_144 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c144
*+ bl_0_144 br_0_144 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c144
*+ bl_0_144 br_0_144 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c144
*+ bl_0_144 br_0_144 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c144
*+ bl_0_144 br_0_144 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c144
*+ bl_0_144 br_0_144 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c144
*+ bl_0_144 br_0_144 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c144
*+ bl_0_144 br_0_144 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c144
*+ bl_0_144 br_0_144 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c144
*+ bl_0_144 br_0_144 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c144
*+ bl_0_144 br_0_144 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c144
*+ bl_0_144 br_0_144 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c144
*+ bl_0_144 br_0_144 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c144
*+ bl_0_144 br_0_144 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c144
*+ bl_0_144 br_0_144 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c144
*+ bl_0_144 br_0_144 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c144
*+ bl_0_144 br_0_144 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c144
*+ bl_0_144 br_0_144 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c144
*+ bl_0_144 br_0_144 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c144
*+ bl_0_144 br_0_144 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c144
*+ bl_0_144 br_0_144 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c144
*+ bl_0_144 br_0_144 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c144
*+ bl_0_144 br_0_144 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c144
*+ bl_0_144 br_0_144 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c144
*+ bl_0_144 br_0_144 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c144
*+ bl_0_144 br_0_144 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c144
*+ bl_0_144 br_0_144 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c144
*+ bl_0_144 br_0_144 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c144
*+ bl_0_144 br_0_144 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c144
*+ bl_0_144 br_0_144 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c144
*+ bl_0_144 br_0_144 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c144
*+ bl_0_144 br_0_144 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c144
*+ bl_0_144 br_0_144 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c144
*+ bl_0_144 br_0_144 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c144
*+ bl_0_144 br_0_144 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c144
*+ bl_0_144 br_0_144 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c144
*+ bl_0_144 br_0_144 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c144
*+ bl_0_144 br_0_144 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c144
*+ bl_0_144 br_0_144 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c144
*+ bl_0_144 br_0_144 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c144
*+ bl_0_144 br_0_144 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c144
*+ bl_0_144 br_0_144 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c144
*+ bl_0_144 br_0_144 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c144
*+ bl_0_144 br_0_144 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c144
*+ bl_0_144 br_0_144 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c144
*+ bl_0_144 br_0_144 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c144
*+ bl_0_144 br_0_144 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c144
*+ bl_0_144 br_0_144 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c144
*+ bl_0_144 br_0_144 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c144
*+ bl_0_144 br_0_144 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c144
*+ bl_0_144 br_0_144 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c144
*+ bl_0_144 br_0_144 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c144
*+ bl_0_144 br_0_144 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c144
*+ bl_0_144 br_0_144 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c144
*+ bl_0_144 br_0_144 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c144
*+ bl_0_144 br_0_144 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c144
*+ bl_0_144 br_0_144 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c144
*+ bl_0_144 br_0_144 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c144
*+ bl_0_144 br_0_144 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c144
*+ bl_0_144 br_0_144 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c144
*+ bl_0_144 br_0_144 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c144
*+ bl_0_144 br_0_144 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c144
*+ bl_0_144 br_0_144 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c144
*+ bl_0_144 br_0_144 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c144
*+ bl_0_144 br_0_144 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c144
*+ bl_0_144 br_0_144 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c144
+ bl_0_144 br_0_144 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c145
+ bl_0_145 br_0_145 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c145
*+ bl_0_145 br_0_145 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c145
*+ bl_0_145 br_0_145 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c145
*+ bl_0_145 br_0_145 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c145
*+ bl_0_145 br_0_145 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c145
*+ bl_0_145 br_0_145 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c145
*+ bl_0_145 br_0_145 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c145
*+ bl_0_145 br_0_145 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c145
*+ bl_0_145 br_0_145 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c145
*+ bl_0_145 br_0_145 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c145
*+ bl_0_145 br_0_145 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c145
*+ bl_0_145 br_0_145 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c145
*+ bl_0_145 br_0_145 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c145
*+ bl_0_145 br_0_145 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c145
*+ bl_0_145 br_0_145 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c145
*+ bl_0_145 br_0_145 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c145
*+ bl_0_145 br_0_145 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c145
*+ bl_0_145 br_0_145 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c145
*+ bl_0_145 br_0_145 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c145
*+ bl_0_145 br_0_145 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c145
*+ bl_0_145 br_0_145 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c145
*+ bl_0_145 br_0_145 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c145
*+ bl_0_145 br_0_145 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c145
*+ bl_0_145 br_0_145 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c145
*+ bl_0_145 br_0_145 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c145
*+ bl_0_145 br_0_145 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c145
*+ bl_0_145 br_0_145 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c145
*+ bl_0_145 br_0_145 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c145
*+ bl_0_145 br_0_145 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c145
*+ bl_0_145 br_0_145 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c145
*+ bl_0_145 br_0_145 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c145
*+ bl_0_145 br_0_145 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c145
*+ bl_0_145 br_0_145 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c145
*+ bl_0_145 br_0_145 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c145
*+ bl_0_145 br_0_145 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c145
*+ bl_0_145 br_0_145 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c145
*+ bl_0_145 br_0_145 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c145
*+ bl_0_145 br_0_145 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c145
*+ bl_0_145 br_0_145 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c145
*+ bl_0_145 br_0_145 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c145
*+ bl_0_145 br_0_145 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c145
*+ bl_0_145 br_0_145 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c145
*+ bl_0_145 br_0_145 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c145
*+ bl_0_145 br_0_145 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c145
*+ bl_0_145 br_0_145 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c145
*+ bl_0_145 br_0_145 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c145
*+ bl_0_145 br_0_145 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c145
*+ bl_0_145 br_0_145 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c145
*+ bl_0_145 br_0_145 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c145
*+ bl_0_145 br_0_145 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c145
*+ bl_0_145 br_0_145 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c145
*+ bl_0_145 br_0_145 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c145
*+ bl_0_145 br_0_145 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c145
*+ bl_0_145 br_0_145 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c145
*+ bl_0_145 br_0_145 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c145
*+ bl_0_145 br_0_145 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c145
*+ bl_0_145 br_0_145 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c145
*+ bl_0_145 br_0_145 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c145
*+ bl_0_145 br_0_145 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c145
*+ bl_0_145 br_0_145 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c145
*+ bl_0_145 br_0_145 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c145
*+ bl_0_145 br_0_145 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c145
*+ bl_0_145 br_0_145 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c145
*+ bl_0_145 br_0_145 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c145
*+ bl_0_145 br_0_145 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c145
*+ bl_0_145 br_0_145 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c145
*+ bl_0_145 br_0_145 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c145
*+ bl_0_145 br_0_145 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c145
*+ bl_0_145 br_0_145 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c145
*+ bl_0_145 br_0_145 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c145
*+ bl_0_145 br_0_145 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c145
*+ bl_0_145 br_0_145 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c145
*+ bl_0_145 br_0_145 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c145
*+ bl_0_145 br_0_145 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c145
*+ bl_0_145 br_0_145 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c145
*+ bl_0_145 br_0_145 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c145
*+ bl_0_145 br_0_145 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c145
*+ bl_0_145 br_0_145 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c145
*+ bl_0_145 br_0_145 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c145
*+ bl_0_145 br_0_145 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c145
*+ bl_0_145 br_0_145 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c145
*+ bl_0_145 br_0_145 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c145
*+ bl_0_145 br_0_145 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c145
*+ bl_0_145 br_0_145 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c145
*+ bl_0_145 br_0_145 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c145
*+ bl_0_145 br_0_145 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c145
*+ bl_0_145 br_0_145 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c145
*+ bl_0_145 br_0_145 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c145
*+ bl_0_145 br_0_145 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c145
*+ bl_0_145 br_0_145 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c145
*+ bl_0_145 br_0_145 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c145
*+ bl_0_145 br_0_145 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c145
*+ bl_0_145 br_0_145 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c145
*+ bl_0_145 br_0_145 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c145
*+ bl_0_145 br_0_145 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c145
*+ bl_0_145 br_0_145 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c145
*+ bl_0_145 br_0_145 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c145
*+ bl_0_145 br_0_145 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c145
*+ bl_0_145 br_0_145 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c145
*+ bl_0_145 br_0_145 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c145
*+ bl_0_145 br_0_145 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c145
*+ bl_0_145 br_0_145 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c145
*+ bl_0_145 br_0_145 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c145
*+ bl_0_145 br_0_145 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c145
*+ bl_0_145 br_0_145 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c145
*+ bl_0_145 br_0_145 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c145
*+ bl_0_145 br_0_145 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c145
*+ bl_0_145 br_0_145 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c145
*+ bl_0_145 br_0_145 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c145
*+ bl_0_145 br_0_145 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c145
*+ bl_0_145 br_0_145 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c145
*+ bl_0_145 br_0_145 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c145
*+ bl_0_145 br_0_145 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c145
*+ bl_0_145 br_0_145 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c145
*+ bl_0_145 br_0_145 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c145
*+ bl_0_145 br_0_145 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c145
*+ bl_0_145 br_0_145 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c145
*+ bl_0_145 br_0_145 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c145
*+ bl_0_145 br_0_145 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c145
*+ bl_0_145 br_0_145 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c145
*+ bl_0_145 br_0_145 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c145
*+ bl_0_145 br_0_145 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c145
*+ bl_0_145 br_0_145 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c145
*+ bl_0_145 br_0_145 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c145
*+ bl_0_145 br_0_145 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c145
*+ bl_0_145 br_0_145 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c145
*+ bl_0_145 br_0_145 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c145
+ bl_0_145 br_0_145 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c146
+ bl_0_146 br_0_146 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c146
*+ bl_0_146 br_0_146 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c146
*+ bl_0_146 br_0_146 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c146
*+ bl_0_146 br_0_146 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c146
*+ bl_0_146 br_0_146 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c146
*+ bl_0_146 br_0_146 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c146
*+ bl_0_146 br_0_146 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c146
*+ bl_0_146 br_0_146 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c146
*+ bl_0_146 br_0_146 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c146
*+ bl_0_146 br_0_146 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c146
*+ bl_0_146 br_0_146 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c146
*+ bl_0_146 br_0_146 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c146
*+ bl_0_146 br_0_146 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c146
*+ bl_0_146 br_0_146 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c146
*+ bl_0_146 br_0_146 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c146
*+ bl_0_146 br_0_146 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c146
*+ bl_0_146 br_0_146 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c146
*+ bl_0_146 br_0_146 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c146
*+ bl_0_146 br_0_146 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c146
*+ bl_0_146 br_0_146 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c146
*+ bl_0_146 br_0_146 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c146
*+ bl_0_146 br_0_146 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c146
*+ bl_0_146 br_0_146 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c146
*+ bl_0_146 br_0_146 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c146
*+ bl_0_146 br_0_146 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c146
*+ bl_0_146 br_0_146 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c146
*+ bl_0_146 br_0_146 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c146
*+ bl_0_146 br_0_146 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c146
*+ bl_0_146 br_0_146 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c146
*+ bl_0_146 br_0_146 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c146
*+ bl_0_146 br_0_146 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c146
*+ bl_0_146 br_0_146 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c146
*+ bl_0_146 br_0_146 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c146
*+ bl_0_146 br_0_146 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c146
*+ bl_0_146 br_0_146 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c146
*+ bl_0_146 br_0_146 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c146
*+ bl_0_146 br_0_146 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c146
*+ bl_0_146 br_0_146 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c146
*+ bl_0_146 br_0_146 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c146
*+ bl_0_146 br_0_146 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c146
*+ bl_0_146 br_0_146 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c146
*+ bl_0_146 br_0_146 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c146
*+ bl_0_146 br_0_146 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c146
*+ bl_0_146 br_0_146 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c146
*+ bl_0_146 br_0_146 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c146
*+ bl_0_146 br_0_146 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c146
*+ bl_0_146 br_0_146 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c146
*+ bl_0_146 br_0_146 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c146
*+ bl_0_146 br_0_146 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c146
*+ bl_0_146 br_0_146 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c146
*+ bl_0_146 br_0_146 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c146
*+ bl_0_146 br_0_146 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c146
*+ bl_0_146 br_0_146 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c146
*+ bl_0_146 br_0_146 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c146
*+ bl_0_146 br_0_146 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c146
*+ bl_0_146 br_0_146 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c146
*+ bl_0_146 br_0_146 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c146
*+ bl_0_146 br_0_146 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c146
*+ bl_0_146 br_0_146 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c146
*+ bl_0_146 br_0_146 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c146
*+ bl_0_146 br_0_146 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c146
*+ bl_0_146 br_0_146 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c146
*+ bl_0_146 br_0_146 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c146
*+ bl_0_146 br_0_146 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c146
*+ bl_0_146 br_0_146 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c146
*+ bl_0_146 br_0_146 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c146
*+ bl_0_146 br_0_146 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c146
*+ bl_0_146 br_0_146 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c146
*+ bl_0_146 br_0_146 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c146
*+ bl_0_146 br_0_146 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c146
*+ bl_0_146 br_0_146 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c146
*+ bl_0_146 br_0_146 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c146
*+ bl_0_146 br_0_146 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c146
*+ bl_0_146 br_0_146 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c146
*+ bl_0_146 br_0_146 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c146
*+ bl_0_146 br_0_146 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c146
*+ bl_0_146 br_0_146 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c146
*+ bl_0_146 br_0_146 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c146
*+ bl_0_146 br_0_146 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c146
*+ bl_0_146 br_0_146 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c146
*+ bl_0_146 br_0_146 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c146
*+ bl_0_146 br_0_146 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c146
*+ bl_0_146 br_0_146 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c146
*+ bl_0_146 br_0_146 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c146
*+ bl_0_146 br_0_146 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c146
*+ bl_0_146 br_0_146 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c146
*+ bl_0_146 br_0_146 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c146
*+ bl_0_146 br_0_146 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c146
*+ bl_0_146 br_0_146 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c146
*+ bl_0_146 br_0_146 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c146
*+ bl_0_146 br_0_146 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c146
*+ bl_0_146 br_0_146 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c146
*+ bl_0_146 br_0_146 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c146
*+ bl_0_146 br_0_146 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c146
*+ bl_0_146 br_0_146 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c146
*+ bl_0_146 br_0_146 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c146
*+ bl_0_146 br_0_146 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c146
*+ bl_0_146 br_0_146 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c146
*+ bl_0_146 br_0_146 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c146
*+ bl_0_146 br_0_146 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c146
*+ bl_0_146 br_0_146 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c146
*+ bl_0_146 br_0_146 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c146
*+ bl_0_146 br_0_146 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c146
*+ bl_0_146 br_0_146 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c146
*+ bl_0_146 br_0_146 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c146
*+ bl_0_146 br_0_146 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c146
*+ bl_0_146 br_0_146 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c146
*+ bl_0_146 br_0_146 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c146
*+ bl_0_146 br_0_146 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c146
*+ bl_0_146 br_0_146 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c146
*+ bl_0_146 br_0_146 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c146
*+ bl_0_146 br_0_146 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c146
*+ bl_0_146 br_0_146 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c146
*+ bl_0_146 br_0_146 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c146
*+ bl_0_146 br_0_146 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c146
*+ bl_0_146 br_0_146 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c146
*+ bl_0_146 br_0_146 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c146
*+ bl_0_146 br_0_146 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c146
*+ bl_0_146 br_0_146 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c146
*+ bl_0_146 br_0_146 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c146
*+ bl_0_146 br_0_146 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c146
*+ bl_0_146 br_0_146 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c146
*+ bl_0_146 br_0_146 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c146
*+ bl_0_146 br_0_146 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c146
*+ bl_0_146 br_0_146 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c146
*+ bl_0_146 br_0_146 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c146
*+ bl_0_146 br_0_146 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c146
+ bl_0_146 br_0_146 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c147
+ bl_0_147 br_0_147 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c147
*+ bl_0_147 br_0_147 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c147
*+ bl_0_147 br_0_147 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c147
*+ bl_0_147 br_0_147 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c147
*+ bl_0_147 br_0_147 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c147
*+ bl_0_147 br_0_147 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c147
*+ bl_0_147 br_0_147 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c147
*+ bl_0_147 br_0_147 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c147
*+ bl_0_147 br_0_147 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c147
*+ bl_0_147 br_0_147 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c147
*+ bl_0_147 br_0_147 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c147
*+ bl_0_147 br_0_147 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c147
*+ bl_0_147 br_0_147 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c147
*+ bl_0_147 br_0_147 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c147
*+ bl_0_147 br_0_147 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c147
*+ bl_0_147 br_0_147 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c147
*+ bl_0_147 br_0_147 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c147
*+ bl_0_147 br_0_147 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c147
*+ bl_0_147 br_0_147 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c147
*+ bl_0_147 br_0_147 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c147
*+ bl_0_147 br_0_147 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c147
*+ bl_0_147 br_0_147 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c147
*+ bl_0_147 br_0_147 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c147
*+ bl_0_147 br_0_147 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c147
*+ bl_0_147 br_0_147 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c147
*+ bl_0_147 br_0_147 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c147
*+ bl_0_147 br_0_147 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c147
*+ bl_0_147 br_0_147 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c147
*+ bl_0_147 br_0_147 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c147
*+ bl_0_147 br_0_147 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c147
*+ bl_0_147 br_0_147 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c147
*+ bl_0_147 br_0_147 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c147
*+ bl_0_147 br_0_147 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c147
*+ bl_0_147 br_0_147 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c147
*+ bl_0_147 br_0_147 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c147
*+ bl_0_147 br_0_147 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c147
*+ bl_0_147 br_0_147 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c147
*+ bl_0_147 br_0_147 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c147
*+ bl_0_147 br_0_147 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c147
*+ bl_0_147 br_0_147 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c147
*+ bl_0_147 br_0_147 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c147
*+ bl_0_147 br_0_147 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c147
*+ bl_0_147 br_0_147 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c147
*+ bl_0_147 br_0_147 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c147
*+ bl_0_147 br_0_147 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c147
*+ bl_0_147 br_0_147 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c147
*+ bl_0_147 br_0_147 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c147
*+ bl_0_147 br_0_147 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c147
*+ bl_0_147 br_0_147 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c147
*+ bl_0_147 br_0_147 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c147
*+ bl_0_147 br_0_147 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c147
*+ bl_0_147 br_0_147 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c147
*+ bl_0_147 br_0_147 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c147
*+ bl_0_147 br_0_147 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c147
*+ bl_0_147 br_0_147 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c147
*+ bl_0_147 br_0_147 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c147
*+ bl_0_147 br_0_147 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c147
*+ bl_0_147 br_0_147 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c147
*+ bl_0_147 br_0_147 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c147
*+ bl_0_147 br_0_147 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c147
*+ bl_0_147 br_0_147 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c147
*+ bl_0_147 br_0_147 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c147
*+ bl_0_147 br_0_147 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c147
*+ bl_0_147 br_0_147 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c147
*+ bl_0_147 br_0_147 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c147
*+ bl_0_147 br_0_147 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c147
*+ bl_0_147 br_0_147 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c147
*+ bl_0_147 br_0_147 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c147
*+ bl_0_147 br_0_147 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c147
*+ bl_0_147 br_0_147 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c147
*+ bl_0_147 br_0_147 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c147
*+ bl_0_147 br_0_147 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c147
*+ bl_0_147 br_0_147 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c147
*+ bl_0_147 br_0_147 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c147
*+ bl_0_147 br_0_147 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c147
*+ bl_0_147 br_0_147 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c147
*+ bl_0_147 br_0_147 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c147
*+ bl_0_147 br_0_147 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c147
*+ bl_0_147 br_0_147 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c147
*+ bl_0_147 br_0_147 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c147
*+ bl_0_147 br_0_147 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c147
*+ bl_0_147 br_0_147 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c147
*+ bl_0_147 br_0_147 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c147
*+ bl_0_147 br_0_147 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c147
*+ bl_0_147 br_0_147 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c147
*+ bl_0_147 br_0_147 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c147
*+ bl_0_147 br_0_147 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c147
*+ bl_0_147 br_0_147 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c147
*+ bl_0_147 br_0_147 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c147
*+ bl_0_147 br_0_147 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c147
*+ bl_0_147 br_0_147 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c147
*+ bl_0_147 br_0_147 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c147
*+ bl_0_147 br_0_147 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c147
*+ bl_0_147 br_0_147 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c147
*+ bl_0_147 br_0_147 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c147
*+ bl_0_147 br_0_147 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c147
*+ bl_0_147 br_0_147 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c147
*+ bl_0_147 br_0_147 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c147
*+ bl_0_147 br_0_147 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c147
*+ bl_0_147 br_0_147 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c147
*+ bl_0_147 br_0_147 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c147
*+ bl_0_147 br_0_147 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c147
*+ bl_0_147 br_0_147 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c147
*+ bl_0_147 br_0_147 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c147
*+ bl_0_147 br_0_147 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c147
*+ bl_0_147 br_0_147 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c147
*+ bl_0_147 br_0_147 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c147
*+ bl_0_147 br_0_147 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c147
*+ bl_0_147 br_0_147 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c147
*+ bl_0_147 br_0_147 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c147
*+ bl_0_147 br_0_147 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c147
*+ bl_0_147 br_0_147 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c147
*+ bl_0_147 br_0_147 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c147
*+ bl_0_147 br_0_147 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c147
*+ bl_0_147 br_0_147 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c147
*+ bl_0_147 br_0_147 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c147
*+ bl_0_147 br_0_147 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c147
*+ bl_0_147 br_0_147 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c147
*+ bl_0_147 br_0_147 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c147
*+ bl_0_147 br_0_147 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c147
*+ bl_0_147 br_0_147 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c147
*+ bl_0_147 br_0_147 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c147
*+ bl_0_147 br_0_147 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c147
*+ bl_0_147 br_0_147 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c147
*+ bl_0_147 br_0_147 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c147
*+ bl_0_147 br_0_147 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c147
*+ bl_0_147 br_0_147 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c147
+ bl_0_147 br_0_147 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c148
+ bl_0_148 br_0_148 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c148
*+ bl_0_148 br_0_148 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c148
*+ bl_0_148 br_0_148 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c148
*+ bl_0_148 br_0_148 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c148
*+ bl_0_148 br_0_148 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c148
*+ bl_0_148 br_0_148 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c148
*+ bl_0_148 br_0_148 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c148
*+ bl_0_148 br_0_148 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c148
*+ bl_0_148 br_0_148 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c148
*+ bl_0_148 br_0_148 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c148
*+ bl_0_148 br_0_148 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c148
*+ bl_0_148 br_0_148 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c148
*+ bl_0_148 br_0_148 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c148
*+ bl_0_148 br_0_148 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c148
*+ bl_0_148 br_0_148 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c148
*+ bl_0_148 br_0_148 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c148
*+ bl_0_148 br_0_148 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c148
*+ bl_0_148 br_0_148 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c148
*+ bl_0_148 br_0_148 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c148
*+ bl_0_148 br_0_148 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c148
*+ bl_0_148 br_0_148 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c148
*+ bl_0_148 br_0_148 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c148
*+ bl_0_148 br_0_148 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c148
*+ bl_0_148 br_0_148 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c148
*+ bl_0_148 br_0_148 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c148
*+ bl_0_148 br_0_148 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c148
*+ bl_0_148 br_0_148 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c148
*+ bl_0_148 br_0_148 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c148
*+ bl_0_148 br_0_148 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c148
*+ bl_0_148 br_0_148 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c148
*+ bl_0_148 br_0_148 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c148
*+ bl_0_148 br_0_148 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c148
*+ bl_0_148 br_0_148 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c148
*+ bl_0_148 br_0_148 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c148
*+ bl_0_148 br_0_148 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c148
*+ bl_0_148 br_0_148 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c148
*+ bl_0_148 br_0_148 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c148
*+ bl_0_148 br_0_148 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c148
*+ bl_0_148 br_0_148 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c148
*+ bl_0_148 br_0_148 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c148
*+ bl_0_148 br_0_148 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c148
*+ bl_0_148 br_0_148 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c148
*+ bl_0_148 br_0_148 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c148
*+ bl_0_148 br_0_148 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c148
*+ bl_0_148 br_0_148 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c148
*+ bl_0_148 br_0_148 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c148
*+ bl_0_148 br_0_148 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c148
*+ bl_0_148 br_0_148 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c148
*+ bl_0_148 br_0_148 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c148
*+ bl_0_148 br_0_148 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c148
*+ bl_0_148 br_0_148 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c148
*+ bl_0_148 br_0_148 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c148
*+ bl_0_148 br_0_148 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c148
*+ bl_0_148 br_0_148 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c148
*+ bl_0_148 br_0_148 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c148
*+ bl_0_148 br_0_148 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c148
*+ bl_0_148 br_0_148 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c148
*+ bl_0_148 br_0_148 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c148
*+ bl_0_148 br_0_148 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c148
*+ bl_0_148 br_0_148 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c148
*+ bl_0_148 br_0_148 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c148
*+ bl_0_148 br_0_148 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c148
*+ bl_0_148 br_0_148 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c148
*+ bl_0_148 br_0_148 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c148
*+ bl_0_148 br_0_148 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c148
*+ bl_0_148 br_0_148 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c148
*+ bl_0_148 br_0_148 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c148
*+ bl_0_148 br_0_148 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c148
*+ bl_0_148 br_0_148 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c148
*+ bl_0_148 br_0_148 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c148
*+ bl_0_148 br_0_148 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c148
*+ bl_0_148 br_0_148 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c148
*+ bl_0_148 br_0_148 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c148
*+ bl_0_148 br_0_148 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c148
*+ bl_0_148 br_0_148 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c148
*+ bl_0_148 br_0_148 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c148
*+ bl_0_148 br_0_148 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c148
*+ bl_0_148 br_0_148 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c148
*+ bl_0_148 br_0_148 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c148
*+ bl_0_148 br_0_148 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c148
*+ bl_0_148 br_0_148 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c148
*+ bl_0_148 br_0_148 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c148
*+ bl_0_148 br_0_148 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c148
*+ bl_0_148 br_0_148 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c148
*+ bl_0_148 br_0_148 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c148
*+ bl_0_148 br_0_148 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c148
*+ bl_0_148 br_0_148 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c148
*+ bl_0_148 br_0_148 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c148
*+ bl_0_148 br_0_148 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c148
*+ bl_0_148 br_0_148 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c148
*+ bl_0_148 br_0_148 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c148
*+ bl_0_148 br_0_148 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c148
*+ bl_0_148 br_0_148 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c148
*+ bl_0_148 br_0_148 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c148
*+ bl_0_148 br_0_148 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c148
*+ bl_0_148 br_0_148 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c148
*+ bl_0_148 br_0_148 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c148
*+ bl_0_148 br_0_148 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c148
*+ bl_0_148 br_0_148 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c148
*+ bl_0_148 br_0_148 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c148
*+ bl_0_148 br_0_148 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c148
*+ bl_0_148 br_0_148 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c148
*+ bl_0_148 br_0_148 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c148
*+ bl_0_148 br_0_148 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c148
*+ bl_0_148 br_0_148 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c148
*+ bl_0_148 br_0_148 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c148
*+ bl_0_148 br_0_148 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c148
*+ bl_0_148 br_0_148 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c148
*+ bl_0_148 br_0_148 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c148
*+ bl_0_148 br_0_148 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c148
*+ bl_0_148 br_0_148 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c148
*+ bl_0_148 br_0_148 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c148
*+ bl_0_148 br_0_148 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c148
*+ bl_0_148 br_0_148 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c148
*+ bl_0_148 br_0_148 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c148
*+ bl_0_148 br_0_148 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c148
*+ bl_0_148 br_0_148 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c148
*+ bl_0_148 br_0_148 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c148
*+ bl_0_148 br_0_148 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c148
*+ bl_0_148 br_0_148 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c148
*+ bl_0_148 br_0_148 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c148
*+ bl_0_148 br_0_148 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c148
*+ bl_0_148 br_0_148 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c148
*+ bl_0_148 br_0_148 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c148
*+ bl_0_148 br_0_148 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c148
*+ bl_0_148 br_0_148 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c148
*+ bl_0_148 br_0_148 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c148
+ bl_0_148 br_0_148 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c149
+ bl_0_149 br_0_149 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c149
*+ bl_0_149 br_0_149 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c149
*+ bl_0_149 br_0_149 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c149
*+ bl_0_149 br_0_149 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c149
*+ bl_0_149 br_0_149 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c149
*+ bl_0_149 br_0_149 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c149
*+ bl_0_149 br_0_149 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c149
*+ bl_0_149 br_0_149 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c149
*+ bl_0_149 br_0_149 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c149
*+ bl_0_149 br_0_149 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c149
*+ bl_0_149 br_0_149 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c149
*+ bl_0_149 br_0_149 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c149
*+ bl_0_149 br_0_149 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c149
*+ bl_0_149 br_0_149 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c149
*+ bl_0_149 br_0_149 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c149
*+ bl_0_149 br_0_149 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c149
*+ bl_0_149 br_0_149 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c149
*+ bl_0_149 br_0_149 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c149
*+ bl_0_149 br_0_149 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c149
*+ bl_0_149 br_0_149 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c149
*+ bl_0_149 br_0_149 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c149
*+ bl_0_149 br_0_149 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c149
*+ bl_0_149 br_0_149 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c149
*+ bl_0_149 br_0_149 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c149
*+ bl_0_149 br_0_149 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c149
*+ bl_0_149 br_0_149 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c149
*+ bl_0_149 br_0_149 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c149
*+ bl_0_149 br_0_149 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c149
*+ bl_0_149 br_0_149 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c149
*+ bl_0_149 br_0_149 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c149
*+ bl_0_149 br_0_149 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c149
*+ bl_0_149 br_0_149 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c149
*+ bl_0_149 br_0_149 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c149
*+ bl_0_149 br_0_149 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c149
*+ bl_0_149 br_0_149 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c149
*+ bl_0_149 br_0_149 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c149
*+ bl_0_149 br_0_149 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c149
*+ bl_0_149 br_0_149 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c149
*+ bl_0_149 br_0_149 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c149
*+ bl_0_149 br_0_149 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c149
*+ bl_0_149 br_0_149 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c149
*+ bl_0_149 br_0_149 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c149
*+ bl_0_149 br_0_149 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c149
*+ bl_0_149 br_0_149 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c149
*+ bl_0_149 br_0_149 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c149
*+ bl_0_149 br_0_149 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c149
*+ bl_0_149 br_0_149 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c149
*+ bl_0_149 br_0_149 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c149
*+ bl_0_149 br_0_149 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c149
*+ bl_0_149 br_0_149 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c149
*+ bl_0_149 br_0_149 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c149
*+ bl_0_149 br_0_149 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c149
*+ bl_0_149 br_0_149 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c149
*+ bl_0_149 br_0_149 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c149
*+ bl_0_149 br_0_149 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c149
*+ bl_0_149 br_0_149 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c149
*+ bl_0_149 br_0_149 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c149
*+ bl_0_149 br_0_149 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c149
*+ bl_0_149 br_0_149 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c149
*+ bl_0_149 br_0_149 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c149
*+ bl_0_149 br_0_149 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c149
*+ bl_0_149 br_0_149 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c149
*+ bl_0_149 br_0_149 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c149
*+ bl_0_149 br_0_149 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c149
*+ bl_0_149 br_0_149 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c149
*+ bl_0_149 br_0_149 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c149
*+ bl_0_149 br_0_149 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c149
*+ bl_0_149 br_0_149 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c149
*+ bl_0_149 br_0_149 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c149
*+ bl_0_149 br_0_149 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c149
*+ bl_0_149 br_0_149 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c149
*+ bl_0_149 br_0_149 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c149
*+ bl_0_149 br_0_149 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c149
*+ bl_0_149 br_0_149 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c149
*+ bl_0_149 br_0_149 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c149
*+ bl_0_149 br_0_149 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c149
*+ bl_0_149 br_0_149 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c149
*+ bl_0_149 br_0_149 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c149
*+ bl_0_149 br_0_149 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c149
*+ bl_0_149 br_0_149 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c149
*+ bl_0_149 br_0_149 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c149
*+ bl_0_149 br_0_149 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c149
*+ bl_0_149 br_0_149 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c149
*+ bl_0_149 br_0_149 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c149
*+ bl_0_149 br_0_149 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c149
*+ bl_0_149 br_0_149 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c149
*+ bl_0_149 br_0_149 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c149
*+ bl_0_149 br_0_149 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c149
*+ bl_0_149 br_0_149 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c149
*+ bl_0_149 br_0_149 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c149
*+ bl_0_149 br_0_149 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c149
*+ bl_0_149 br_0_149 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c149
*+ bl_0_149 br_0_149 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c149
*+ bl_0_149 br_0_149 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c149
*+ bl_0_149 br_0_149 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c149
*+ bl_0_149 br_0_149 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c149
*+ bl_0_149 br_0_149 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c149
*+ bl_0_149 br_0_149 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c149
*+ bl_0_149 br_0_149 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c149
*+ bl_0_149 br_0_149 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c149
*+ bl_0_149 br_0_149 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c149
*+ bl_0_149 br_0_149 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c149
*+ bl_0_149 br_0_149 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c149
*+ bl_0_149 br_0_149 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c149
*+ bl_0_149 br_0_149 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c149
*+ bl_0_149 br_0_149 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c149
*+ bl_0_149 br_0_149 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c149
*+ bl_0_149 br_0_149 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c149
*+ bl_0_149 br_0_149 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c149
*+ bl_0_149 br_0_149 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c149
*+ bl_0_149 br_0_149 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c149
*+ bl_0_149 br_0_149 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c149
*+ bl_0_149 br_0_149 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c149
*+ bl_0_149 br_0_149 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c149
*+ bl_0_149 br_0_149 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c149
*+ bl_0_149 br_0_149 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c149
*+ bl_0_149 br_0_149 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c149
*+ bl_0_149 br_0_149 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c149
*+ bl_0_149 br_0_149 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c149
*+ bl_0_149 br_0_149 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c149
*+ bl_0_149 br_0_149 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c149
*+ bl_0_149 br_0_149 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c149
*+ bl_0_149 br_0_149 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c149
*+ bl_0_149 br_0_149 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c149
*+ bl_0_149 br_0_149 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c149
*+ bl_0_149 br_0_149 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c149
*+ bl_0_149 br_0_149 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c149
+ bl_0_149 br_0_149 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c150
+ bl_0_150 br_0_150 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c150
*+ bl_0_150 br_0_150 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c150
*+ bl_0_150 br_0_150 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c150
*+ bl_0_150 br_0_150 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c150
*+ bl_0_150 br_0_150 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c150
*+ bl_0_150 br_0_150 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c150
*+ bl_0_150 br_0_150 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c150
*+ bl_0_150 br_0_150 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c150
*+ bl_0_150 br_0_150 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c150
*+ bl_0_150 br_0_150 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c150
*+ bl_0_150 br_0_150 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c150
*+ bl_0_150 br_0_150 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c150
*+ bl_0_150 br_0_150 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c150
*+ bl_0_150 br_0_150 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c150
*+ bl_0_150 br_0_150 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c150
*+ bl_0_150 br_0_150 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c150
*+ bl_0_150 br_0_150 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c150
*+ bl_0_150 br_0_150 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c150
*+ bl_0_150 br_0_150 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c150
*+ bl_0_150 br_0_150 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c150
*+ bl_0_150 br_0_150 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c150
*+ bl_0_150 br_0_150 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c150
*+ bl_0_150 br_0_150 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c150
*+ bl_0_150 br_0_150 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c150
*+ bl_0_150 br_0_150 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c150
*+ bl_0_150 br_0_150 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c150
*+ bl_0_150 br_0_150 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c150
*+ bl_0_150 br_0_150 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c150
*+ bl_0_150 br_0_150 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c150
*+ bl_0_150 br_0_150 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c150
*+ bl_0_150 br_0_150 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c150
*+ bl_0_150 br_0_150 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c150
*+ bl_0_150 br_0_150 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c150
*+ bl_0_150 br_0_150 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c150
*+ bl_0_150 br_0_150 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c150
*+ bl_0_150 br_0_150 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c150
*+ bl_0_150 br_0_150 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c150
*+ bl_0_150 br_0_150 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c150
*+ bl_0_150 br_0_150 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c150
*+ bl_0_150 br_0_150 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c150
*+ bl_0_150 br_0_150 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c150
*+ bl_0_150 br_0_150 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c150
*+ bl_0_150 br_0_150 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c150
*+ bl_0_150 br_0_150 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c150
*+ bl_0_150 br_0_150 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c150
*+ bl_0_150 br_0_150 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c150
*+ bl_0_150 br_0_150 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c150
*+ bl_0_150 br_0_150 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c150
*+ bl_0_150 br_0_150 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c150
*+ bl_0_150 br_0_150 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c150
*+ bl_0_150 br_0_150 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c150
*+ bl_0_150 br_0_150 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c150
*+ bl_0_150 br_0_150 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c150
*+ bl_0_150 br_0_150 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c150
*+ bl_0_150 br_0_150 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c150
*+ bl_0_150 br_0_150 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c150
*+ bl_0_150 br_0_150 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c150
*+ bl_0_150 br_0_150 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c150
*+ bl_0_150 br_0_150 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c150
*+ bl_0_150 br_0_150 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c150
*+ bl_0_150 br_0_150 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c150
*+ bl_0_150 br_0_150 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c150
*+ bl_0_150 br_0_150 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c150
*+ bl_0_150 br_0_150 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c150
*+ bl_0_150 br_0_150 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c150
*+ bl_0_150 br_0_150 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c150
*+ bl_0_150 br_0_150 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c150
*+ bl_0_150 br_0_150 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c150
*+ bl_0_150 br_0_150 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c150
*+ bl_0_150 br_0_150 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c150
*+ bl_0_150 br_0_150 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c150
*+ bl_0_150 br_0_150 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c150
*+ bl_0_150 br_0_150 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c150
*+ bl_0_150 br_0_150 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c150
*+ bl_0_150 br_0_150 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c150
*+ bl_0_150 br_0_150 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c150
*+ bl_0_150 br_0_150 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c150
*+ bl_0_150 br_0_150 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c150
*+ bl_0_150 br_0_150 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c150
*+ bl_0_150 br_0_150 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c150
*+ bl_0_150 br_0_150 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c150
*+ bl_0_150 br_0_150 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c150
*+ bl_0_150 br_0_150 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c150
*+ bl_0_150 br_0_150 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c150
*+ bl_0_150 br_0_150 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c150
*+ bl_0_150 br_0_150 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c150
*+ bl_0_150 br_0_150 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c150
*+ bl_0_150 br_0_150 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c150
*+ bl_0_150 br_0_150 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c150
*+ bl_0_150 br_0_150 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c150
*+ bl_0_150 br_0_150 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c150
*+ bl_0_150 br_0_150 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c150
*+ bl_0_150 br_0_150 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c150
*+ bl_0_150 br_0_150 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c150
*+ bl_0_150 br_0_150 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c150
*+ bl_0_150 br_0_150 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c150
*+ bl_0_150 br_0_150 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c150
*+ bl_0_150 br_0_150 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c150
*+ bl_0_150 br_0_150 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c150
*+ bl_0_150 br_0_150 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c150
*+ bl_0_150 br_0_150 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c150
*+ bl_0_150 br_0_150 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c150
*+ bl_0_150 br_0_150 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c150
*+ bl_0_150 br_0_150 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c150
*+ bl_0_150 br_0_150 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c150
*+ bl_0_150 br_0_150 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c150
*+ bl_0_150 br_0_150 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c150
*+ bl_0_150 br_0_150 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c150
*+ bl_0_150 br_0_150 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c150
*+ bl_0_150 br_0_150 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c150
*+ bl_0_150 br_0_150 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c150
*+ bl_0_150 br_0_150 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c150
*+ bl_0_150 br_0_150 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c150
*+ bl_0_150 br_0_150 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c150
*+ bl_0_150 br_0_150 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c150
*+ bl_0_150 br_0_150 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c150
*+ bl_0_150 br_0_150 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c150
*+ bl_0_150 br_0_150 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c150
*+ bl_0_150 br_0_150 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c150
*+ bl_0_150 br_0_150 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c150
*+ bl_0_150 br_0_150 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c150
*+ bl_0_150 br_0_150 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c150
*+ bl_0_150 br_0_150 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c150
*+ bl_0_150 br_0_150 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c150
*+ bl_0_150 br_0_150 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c150
*+ bl_0_150 br_0_150 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c150
*+ bl_0_150 br_0_150 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c150
+ bl_0_150 br_0_150 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c151
+ bl_0_151 br_0_151 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c151
*+ bl_0_151 br_0_151 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c151
*+ bl_0_151 br_0_151 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c151
*+ bl_0_151 br_0_151 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c151
*+ bl_0_151 br_0_151 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c151
*+ bl_0_151 br_0_151 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c151
*+ bl_0_151 br_0_151 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c151
*+ bl_0_151 br_0_151 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c151
*+ bl_0_151 br_0_151 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c151
*+ bl_0_151 br_0_151 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c151
*+ bl_0_151 br_0_151 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c151
*+ bl_0_151 br_0_151 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c151
*+ bl_0_151 br_0_151 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c151
*+ bl_0_151 br_0_151 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c151
*+ bl_0_151 br_0_151 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c151
*+ bl_0_151 br_0_151 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c151
*+ bl_0_151 br_0_151 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c151
*+ bl_0_151 br_0_151 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c151
*+ bl_0_151 br_0_151 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c151
*+ bl_0_151 br_0_151 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c151
*+ bl_0_151 br_0_151 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c151
*+ bl_0_151 br_0_151 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c151
*+ bl_0_151 br_0_151 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c151
*+ bl_0_151 br_0_151 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c151
*+ bl_0_151 br_0_151 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c151
*+ bl_0_151 br_0_151 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c151
*+ bl_0_151 br_0_151 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c151
*+ bl_0_151 br_0_151 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c151
*+ bl_0_151 br_0_151 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c151
*+ bl_0_151 br_0_151 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c151
*+ bl_0_151 br_0_151 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c151
*+ bl_0_151 br_0_151 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c151
*+ bl_0_151 br_0_151 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c151
*+ bl_0_151 br_0_151 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c151
*+ bl_0_151 br_0_151 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c151
*+ bl_0_151 br_0_151 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c151
*+ bl_0_151 br_0_151 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c151
*+ bl_0_151 br_0_151 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c151
*+ bl_0_151 br_0_151 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c151
*+ bl_0_151 br_0_151 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c151
*+ bl_0_151 br_0_151 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c151
*+ bl_0_151 br_0_151 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c151
*+ bl_0_151 br_0_151 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c151
*+ bl_0_151 br_0_151 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c151
*+ bl_0_151 br_0_151 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c151
*+ bl_0_151 br_0_151 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c151
*+ bl_0_151 br_0_151 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c151
*+ bl_0_151 br_0_151 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c151
*+ bl_0_151 br_0_151 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c151
*+ bl_0_151 br_0_151 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c151
*+ bl_0_151 br_0_151 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c151
*+ bl_0_151 br_0_151 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c151
*+ bl_0_151 br_0_151 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c151
*+ bl_0_151 br_0_151 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c151
*+ bl_0_151 br_0_151 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c151
*+ bl_0_151 br_0_151 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c151
*+ bl_0_151 br_0_151 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c151
*+ bl_0_151 br_0_151 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c151
*+ bl_0_151 br_0_151 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c151
*+ bl_0_151 br_0_151 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c151
*+ bl_0_151 br_0_151 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c151
*+ bl_0_151 br_0_151 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c151
*+ bl_0_151 br_0_151 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c151
*+ bl_0_151 br_0_151 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c151
*+ bl_0_151 br_0_151 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c151
*+ bl_0_151 br_0_151 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c151
*+ bl_0_151 br_0_151 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c151
*+ bl_0_151 br_0_151 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c151
*+ bl_0_151 br_0_151 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c151
*+ bl_0_151 br_0_151 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c151
*+ bl_0_151 br_0_151 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c151
*+ bl_0_151 br_0_151 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c151
*+ bl_0_151 br_0_151 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c151
*+ bl_0_151 br_0_151 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c151
*+ bl_0_151 br_0_151 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c151
*+ bl_0_151 br_0_151 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c151
*+ bl_0_151 br_0_151 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c151
*+ bl_0_151 br_0_151 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c151
*+ bl_0_151 br_0_151 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c151
*+ bl_0_151 br_0_151 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c151
*+ bl_0_151 br_0_151 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c151
*+ bl_0_151 br_0_151 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c151
*+ bl_0_151 br_0_151 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c151
*+ bl_0_151 br_0_151 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c151
*+ bl_0_151 br_0_151 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c151
*+ bl_0_151 br_0_151 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c151
*+ bl_0_151 br_0_151 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c151
*+ bl_0_151 br_0_151 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c151
*+ bl_0_151 br_0_151 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c151
*+ bl_0_151 br_0_151 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c151
*+ bl_0_151 br_0_151 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c151
*+ bl_0_151 br_0_151 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c151
*+ bl_0_151 br_0_151 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c151
*+ bl_0_151 br_0_151 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c151
*+ bl_0_151 br_0_151 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c151
*+ bl_0_151 br_0_151 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c151
*+ bl_0_151 br_0_151 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c151
*+ bl_0_151 br_0_151 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c151
*+ bl_0_151 br_0_151 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c151
*+ bl_0_151 br_0_151 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c151
*+ bl_0_151 br_0_151 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c151
*+ bl_0_151 br_0_151 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c151
*+ bl_0_151 br_0_151 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c151
*+ bl_0_151 br_0_151 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c151
*+ bl_0_151 br_0_151 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c151
*+ bl_0_151 br_0_151 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c151
*+ bl_0_151 br_0_151 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c151
*+ bl_0_151 br_0_151 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c151
*+ bl_0_151 br_0_151 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c151
*+ bl_0_151 br_0_151 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c151
*+ bl_0_151 br_0_151 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c151
*+ bl_0_151 br_0_151 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c151
*+ bl_0_151 br_0_151 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c151
*+ bl_0_151 br_0_151 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c151
*+ bl_0_151 br_0_151 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c151
*+ bl_0_151 br_0_151 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c151
*+ bl_0_151 br_0_151 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c151
*+ bl_0_151 br_0_151 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c151
*+ bl_0_151 br_0_151 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c151
*+ bl_0_151 br_0_151 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c151
*+ bl_0_151 br_0_151 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c151
*+ bl_0_151 br_0_151 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c151
*+ bl_0_151 br_0_151 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c151
*+ bl_0_151 br_0_151 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c151
*+ bl_0_151 br_0_151 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c151
*+ bl_0_151 br_0_151 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c151
*+ bl_0_151 br_0_151 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c151
+ bl_0_151 br_0_151 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c152
+ bl_0_152 br_0_152 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c152
*+ bl_0_152 br_0_152 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c152
*+ bl_0_152 br_0_152 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c152
*+ bl_0_152 br_0_152 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c152
*+ bl_0_152 br_0_152 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c152
*+ bl_0_152 br_0_152 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c152
*+ bl_0_152 br_0_152 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c152
*+ bl_0_152 br_0_152 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c152
*+ bl_0_152 br_0_152 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c152
*+ bl_0_152 br_0_152 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c152
*+ bl_0_152 br_0_152 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c152
*+ bl_0_152 br_0_152 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c152
*+ bl_0_152 br_0_152 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c152
*+ bl_0_152 br_0_152 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c152
*+ bl_0_152 br_0_152 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c152
*+ bl_0_152 br_0_152 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c152
*+ bl_0_152 br_0_152 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c152
*+ bl_0_152 br_0_152 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c152
*+ bl_0_152 br_0_152 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c152
*+ bl_0_152 br_0_152 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c152
*+ bl_0_152 br_0_152 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c152
*+ bl_0_152 br_0_152 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c152
*+ bl_0_152 br_0_152 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c152
*+ bl_0_152 br_0_152 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c152
*+ bl_0_152 br_0_152 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c152
*+ bl_0_152 br_0_152 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c152
*+ bl_0_152 br_0_152 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c152
*+ bl_0_152 br_0_152 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c152
*+ bl_0_152 br_0_152 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c152
*+ bl_0_152 br_0_152 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c152
*+ bl_0_152 br_0_152 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c152
*+ bl_0_152 br_0_152 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c152
*+ bl_0_152 br_0_152 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c152
*+ bl_0_152 br_0_152 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c152
*+ bl_0_152 br_0_152 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c152
*+ bl_0_152 br_0_152 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c152
*+ bl_0_152 br_0_152 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c152
*+ bl_0_152 br_0_152 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c152
*+ bl_0_152 br_0_152 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c152
*+ bl_0_152 br_0_152 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c152
*+ bl_0_152 br_0_152 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c152
*+ bl_0_152 br_0_152 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c152
*+ bl_0_152 br_0_152 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c152
*+ bl_0_152 br_0_152 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c152
*+ bl_0_152 br_0_152 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c152
*+ bl_0_152 br_0_152 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c152
*+ bl_0_152 br_0_152 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c152
*+ bl_0_152 br_0_152 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c152
*+ bl_0_152 br_0_152 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c152
*+ bl_0_152 br_0_152 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c152
*+ bl_0_152 br_0_152 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c152
*+ bl_0_152 br_0_152 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c152
*+ bl_0_152 br_0_152 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c152
*+ bl_0_152 br_0_152 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c152
*+ bl_0_152 br_0_152 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c152
*+ bl_0_152 br_0_152 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c152
*+ bl_0_152 br_0_152 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c152
*+ bl_0_152 br_0_152 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c152
*+ bl_0_152 br_0_152 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c152
*+ bl_0_152 br_0_152 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c152
*+ bl_0_152 br_0_152 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c152
*+ bl_0_152 br_0_152 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c152
*+ bl_0_152 br_0_152 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c152
*+ bl_0_152 br_0_152 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c152
*+ bl_0_152 br_0_152 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c152
*+ bl_0_152 br_0_152 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c152
*+ bl_0_152 br_0_152 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c152
*+ bl_0_152 br_0_152 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c152
*+ bl_0_152 br_0_152 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c152
*+ bl_0_152 br_0_152 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c152
*+ bl_0_152 br_0_152 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c152
*+ bl_0_152 br_0_152 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c152
*+ bl_0_152 br_0_152 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c152
*+ bl_0_152 br_0_152 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c152
*+ bl_0_152 br_0_152 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c152
*+ bl_0_152 br_0_152 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c152
*+ bl_0_152 br_0_152 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c152
*+ bl_0_152 br_0_152 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c152
*+ bl_0_152 br_0_152 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c152
*+ bl_0_152 br_0_152 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c152
*+ bl_0_152 br_0_152 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c152
*+ bl_0_152 br_0_152 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c152
*+ bl_0_152 br_0_152 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c152
*+ bl_0_152 br_0_152 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c152
*+ bl_0_152 br_0_152 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c152
*+ bl_0_152 br_0_152 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c152
*+ bl_0_152 br_0_152 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c152
*+ bl_0_152 br_0_152 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c152
*+ bl_0_152 br_0_152 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c152
*+ bl_0_152 br_0_152 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c152
*+ bl_0_152 br_0_152 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c152
*+ bl_0_152 br_0_152 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c152
*+ bl_0_152 br_0_152 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c152
*+ bl_0_152 br_0_152 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c152
*+ bl_0_152 br_0_152 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c152
*+ bl_0_152 br_0_152 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c152
*+ bl_0_152 br_0_152 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c152
*+ bl_0_152 br_0_152 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c152
*+ bl_0_152 br_0_152 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c152
*+ bl_0_152 br_0_152 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c152
*+ bl_0_152 br_0_152 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c152
*+ bl_0_152 br_0_152 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c152
*+ bl_0_152 br_0_152 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c152
*+ bl_0_152 br_0_152 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c152
*+ bl_0_152 br_0_152 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c152
*+ bl_0_152 br_0_152 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c152
*+ bl_0_152 br_0_152 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c152
*+ bl_0_152 br_0_152 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c152
*+ bl_0_152 br_0_152 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c152
*+ bl_0_152 br_0_152 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c152
*+ bl_0_152 br_0_152 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c152
*+ bl_0_152 br_0_152 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c152
*+ bl_0_152 br_0_152 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c152
*+ bl_0_152 br_0_152 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c152
*+ bl_0_152 br_0_152 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c152
*+ bl_0_152 br_0_152 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c152
*+ bl_0_152 br_0_152 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c152
*+ bl_0_152 br_0_152 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c152
*+ bl_0_152 br_0_152 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c152
*+ bl_0_152 br_0_152 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c152
*+ bl_0_152 br_0_152 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c152
*+ bl_0_152 br_0_152 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c152
*+ bl_0_152 br_0_152 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c152
*+ bl_0_152 br_0_152 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c152
*+ bl_0_152 br_0_152 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c152
*+ bl_0_152 br_0_152 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c152
*+ bl_0_152 br_0_152 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c152
+ bl_0_152 br_0_152 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c153
+ bl_0_153 br_0_153 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c153
*+ bl_0_153 br_0_153 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c153
*+ bl_0_153 br_0_153 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c153
*+ bl_0_153 br_0_153 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c153
*+ bl_0_153 br_0_153 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c153
*+ bl_0_153 br_0_153 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c153
*+ bl_0_153 br_0_153 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c153
*+ bl_0_153 br_0_153 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c153
*+ bl_0_153 br_0_153 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c153
*+ bl_0_153 br_0_153 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c153
*+ bl_0_153 br_0_153 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c153
*+ bl_0_153 br_0_153 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c153
*+ bl_0_153 br_0_153 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c153
*+ bl_0_153 br_0_153 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c153
*+ bl_0_153 br_0_153 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c153
*+ bl_0_153 br_0_153 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c153
*+ bl_0_153 br_0_153 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c153
*+ bl_0_153 br_0_153 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c153
*+ bl_0_153 br_0_153 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c153
*+ bl_0_153 br_0_153 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c153
*+ bl_0_153 br_0_153 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c153
*+ bl_0_153 br_0_153 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c153
*+ bl_0_153 br_0_153 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c153
*+ bl_0_153 br_0_153 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c153
*+ bl_0_153 br_0_153 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c153
*+ bl_0_153 br_0_153 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c153
*+ bl_0_153 br_0_153 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c153
*+ bl_0_153 br_0_153 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c153
*+ bl_0_153 br_0_153 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c153
*+ bl_0_153 br_0_153 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c153
*+ bl_0_153 br_0_153 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c153
*+ bl_0_153 br_0_153 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c153
*+ bl_0_153 br_0_153 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c153
*+ bl_0_153 br_0_153 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c153
*+ bl_0_153 br_0_153 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c153
*+ bl_0_153 br_0_153 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c153
*+ bl_0_153 br_0_153 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c153
*+ bl_0_153 br_0_153 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c153
*+ bl_0_153 br_0_153 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c153
*+ bl_0_153 br_0_153 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c153
*+ bl_0_153 br_0_153 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c153
*+ bl_0_153 br_0_153 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c153
*+ bl_0_153 br_0_153 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c153
*+ bl_0_153 br_0_153 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c153
*+ bl_0_153 br_0_153 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c153
*+ bl_0_153 br_0_153 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c153
*+ bl_0_153 br_0_153 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c153
*+ bl_0_153 br_0_153 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c153
*+ bl_0_153 br_0_153 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c153
*+ bl_0_153 br_0_153 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c153
*+ bl_0_153 br_0_153 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c153
*+ bl_0_153 br_0_153 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c153
*+ bl_0_153 br_0_153 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c153
*+ bl_0_153 br_0_153 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c153
*+ bl_0_153 br_0_153 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c153
*+ bl_0_153 br_0_153 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c153
*+ bl_0_153 br_0_153 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c153
*+ bl_0_153 br_0_153 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c153
*+ bl_0_153 br_0_153 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c153
*+ bl_0_153 br_0_153 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c153
*+ bl_0_153 br_0_153 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c153
*+ bl_0_153 br_0_153 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c153
*+ bl_0_153 br_0_153 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c153
*+ bl_0_153 br_0_153 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c153
*+ bl_0_153 br_0_153 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c153
*+ bl_0_153 br_0_153 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c153
*+ bl_0_153 br_0_153 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c153
*+ bl_0_153 br_0_153 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c153
*+ bl_0_153 br_0_153 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c153
*+ bl_0_153 br_0_153 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c153
*+ bl_0_153 br_0_153 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c153
*+ bl_0_153 br_0_153 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c153
*+ bl_0_153 br_0_153 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c153
*+ bl_0_153 br_0_153 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c153
*+ bl_0_153 br_0_153 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c153
*+ bl_0_153 br_0_153 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c153
*+ bl_0_153 br_0_153 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c153
*+ bl_0_153 br_0_153 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c153
*+ bl_0_153 br_0_153 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c153
*+ bl_0_153 br_0_153 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c153
*+ bl_0_153 br_0_153 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c153
*+ bl_0_153 br_0_153 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c153
*+ bl_0_153 br_0_153 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c153
*+ bl_0_153 br_0_153 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c153
*+ bl_0_153 br_0_153 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c153
*+ bl_0_153 br_0_153 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c153
*+ bl_0_153 br_0_153 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c153
*+ bl_0_153 br_0_153 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c153
*+ bl_0_153 br_0_153 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c153
*+ bl_0_153 br_0_153 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c153
*+ bl_0_153 br_0_153 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c153
*+ bl_0_153 br_0_153 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c153
*+ bl_0_153 br_0_153 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c153
*+ bl_0_153 br_0_153 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c153
*+ bl_0_153 br_0_153 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c153
*+ bl_0_153 br_0_153 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c153
*+ bl_0_153 br_0_153 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c153
*+ bl_0_153 br_0_153 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c153
*+ bl_0_153 br_0_153 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c153
*+ bl_0_153 br_0_153 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c153
*+ bl_0_153 br_0_153 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c153
*+ bl_0_153 br_0_153 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c153
*+ bl_0_153 br_0_153 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c153
*+ bl_0_153 br_0_153 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c153
*+ bl_0_153 br_0_153 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c153
*+ bl_0_153 br_0_153 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c153
*+ bl_0_153 br_0_153 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c153
*+ bl_0_153 br_0_153 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c153
*+ bl_0_153 br_0_153 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c153
*+ bl_0_153 br_0_153 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c153
*+ bl_0_153 br_0_153 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c153
*+ bl_0_153 br_0_153 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c153
*+ bl_0_153 br_0_153 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c153
*+ bl_0_153 br_0_153 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c153
*+ bl_0_153 br_0_153 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c153
*+ bl_0_153 br_0_153 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c153
*+ bl_0_153 br_0_153 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c153
*+ bl_0_153 br_0_153 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c153
*+ bl_0_153 br_0_153 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c153
*+ bl_0_153 br_0_153 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c153
*+ bl_0_153 br_0_153 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c153
*+ bl_0_153 br_0_153 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c153
*+ bl_0_153 br_0_153 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c153
*+ bl_0_153 br_0_153 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c153
*+ bl_0_153 br_0_153 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c153
*+ bl_0_153 br_0_153 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c153
*+ bl_0_153 br_0_153 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c153
+ bl_0_153 br_0_153 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c154
+ bl_0_154 br_0_154 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c154
*+ bl_0_154 br_0_154 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c154
*+ bl_0_154 br_0_154 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c154
*+ bl_0_154 br_0_154 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c154
*+ bl_0_154 br_0_154 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c154
*+ bl_0_154 br_0_154 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c154
*+ bl_0_154 br_0_154 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c154
*+ bl_0_154 br_0_154 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c154
*+ bl_0_154 br_0_154 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c154
*+ bl_0_154 br_0_154 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c154
*+ bl_0_154 br_0_154 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c154
*+ bl_0_154 br_0_154 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c154
*+ bl_0_154 br_0_154 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c154
*+ bl_0_154 br_0_154 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c154
*+ bl_0_154 br_0_154 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c154
*+ bl_0_154 br_0_154 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c154
*+ bl_0_154 br_0_154 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c154
*+ bl_0_154 br_0_154 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c154
*+ bl_0_154 br_0_154 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c154
*+ bl_0_154 br_0_154 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c154
*+ bl_0_154 br_0_154 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c154
*+ bl_0_154 br_0_154 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c154
*+ bl_0_154 br_0_154 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c154
*+ bl_0_154 br_0_154 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c154
*+ bl_0_154 br_0_154 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c154
*+ bl_0_154 br_0_154 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c154
*+ bl_0_154 br_0_154 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c154
*+ bl_0_154 br_0_154 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c154
*+ bl_0_154 br_0_154 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c154
*+ bl_0_154 br_0_154 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c154
*+ bl_0_154 br_0_154 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c154
*+ bl_0_154 br_0_154 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c154
*+ bl_0_154 br_0_154 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c154
*+ bl_0_154 br_0_154 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c154
*+ bl_0_154 br_0_154 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c154
*+ bl_0_154 br_0_154 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c154
*+ bl_0_154 br_0_154 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c154
*+ bl_0_154 br_0_154 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c154
*+ bl_0_154 br_0_154 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c154
*+ bl_0_154 br_0_154 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c154
*+ bl_0_154 br_0_154 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c154
*+ bl_0_154 br_0_154 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c154
*+ bl_0_154 br_0_154 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c154
*+ bl_0_154 br_0_154 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c154
*+ bl_0_154 br_0_154 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c154
*+ bl_0_154 br_0_154 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c154
*+ bl_0_154 br_0_154 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c154
*+ bl_0_154 br_0_154 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c154
*+ bl_0_154 br_0_154 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c154
*+ bl_0_154 br_0_154 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c154
*+ bl_0_154 br_0_154 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c154
*+ bl_0_154 br_0_154 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c154
*+ bl_0_154 br_0_154 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c154
*+ bl_0_154 br_0_154 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c154
*+ bl_0_154 br_0_154 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c154
*+ bl_0_154 br_0_154 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c154
*+ bl_0_154 br_0_154 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c154
*+ bl_0_154 br_0_154 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c154
*+ bl_0_154 br_0_154 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c154
*+ bl_0_154 br_0_154 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c154
*+ bl_0_154 br_0_154 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c154
*+ bl_0_154 br_0_154 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c154
*+ bl_0_154 br_0_154 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c154
*+ bl_0_154 br_0_154 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c154
*+ bl_0_154 br_0_154 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c154
*+ bl_0_154 br_0_154 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c154
*+ bl_0_154 br_0_154 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c154
*+ bl_0_154 br_0_154 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c154
*+ bl_0_154 br_0_154 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c154
*+ bl_0_154 br_0_154 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c154
*+ bl_0_154 br_0_154 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c154
*+ bl_0_154 br_0_154 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c154
*+ bl_0_154 br_0_154 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c154
*+ bl_0_154 br_0_154 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c154
*+ bl_0_154 br_0_154 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c154
*+ bl_0_154 br_0_154 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c154
*+ bl_0_154 br_0_154 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c154
*+ bl_0_154 br_0_154 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c154
*+ bl_0_154 br_0_154 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c154
*+ bl_0_154 br_0_154 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c154
*+ bl_0_154 br_0_154 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c154
*+ bl_0_154 br_0_154 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c154
*+ bl_0_154 br_0_154 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c154
*+ bl_0_154 br_0_154 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c154
*+ bl_0_154 br_0_154 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c154
*+ bl_0_154 br_0_154 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c154
*+ bl_0_154 br_0_154 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c154
*+ bl_0_154 br_0_154 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c154
*+ bl_0_154 br_0_154 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c154
*+ bl_0_154 br_0_154 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c154
*+ bl_0_154 br_0_154 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c154
*+ bl_0_154 br_0_154 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c154
*+ bl_0_154 br_0_154 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c154
*+ bl_0_154 br_0_154 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c154
*+ bl_0_154 br_0_154 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c154
*+ bl_0_154 br_0_154 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c154
*+ bl_0_154 br_0_154 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c154
*+ bl_0_154 br_0_154 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c154
*+ bl_0_154 br_0_154 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c154
*+ bl_0_154 br_0_154 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c154
*+ bl_0_154 br_0_154 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c154
*+ bl_0_154 br_0_154 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c154
*+ bl_0_154 br_0_154 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c154
*+ bl_0_154 br_0_154 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c154
*+ bl_0_154 br_0_154 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c154
*+ bl_0_154 br_0_154 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c154
*+ bl_0_154 br_0_154 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c154
*+ bl_0_154 br_0_154 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c154
*+ bl_0_154 br_0_154 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c154
*+ bl_0_154 br_0_154 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c154
*+ bl_0_154 br_0_154 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c154
*+ bl_0_154 br_0_154 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c154
*+ bl_0_154 br_0_154 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c154
*+ bl_0_154 br_0_154 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c154
*+ bl_0_154 br_0_154 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c154
*+ bl_0_154 br_0_154 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c154
*+ bl_0_154 br_0_154 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c154
*+ bl_0_154 br_0_154 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c154
*+ bl_0_154 br_0_154 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c154
*+ bl_0_154 br_0_154 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c154
*+ bl_0_154 br_0_154 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c154
*+ bl_0_154 br_0_154 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c154
*+ bl_0_154 br_0_154 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c154
*+ bl_0_154 br_0_154 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c154
*+ bl_0_154 br_0_154 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c154
*+ bl_0_154 br_0_154 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c154
*+ bl_0_154 br_0_154 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c154
+ bl_0_154 br_0_154 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c155
+ bl_0_155 br_0_155 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c155
*+ bl_0_155 br_0_155 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c155
*+ bl_0_155 br_0_155 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c155
*+ bl_0_155 br_0_155 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c155
*+ bl_0_155 br_0_155 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c155
*+ bl_0_155 br_0_155 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c155
*+ bl_0_155 br_0_155 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c155
*+ bl_0_155 br_0_155 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c155
*+ bl_0_155 br_0_155 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c155
*+ bl_0_155 br_0_155 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c155
*+ bl_0_155 br_0_155 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c155
*+ bl_0_155 br_0_155 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c155
*+ bl_0_155 br_0_155 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c155
*+ bl_0_155 br_0_155 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c155
*+ bl_0_155 br_0_155 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c155
*+ bl_0_155 br_0_155 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c155
*+ bl_0_155 br_0_155 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c155
*+ bl_0_155 br_0_155 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c155
*+ bl_0_155 br_0_155 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c155
*+ bl_0_155 br_0_155 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c155
*+ bl_0_155 br_0_155 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c155
*+ bl_0_155 br_0_155 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c155
*+ bl_0_155 br_0_155 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c155
*+ bl_0_155 br_0_155 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c155
*+ bl_0_155 br_0_155 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c155
*+ bl_0_155 br_0_155 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c155
*+ bl_0_155 br_0_155 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c155
*+ bl_0_155 br_0_155 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c155
*+ bl_0_155 br_0_155 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c155
*+ bl_0_155 br_0_155 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c155
*+ bl_0_155 br_0_155 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c155
*+ bl_0_155 br_0_155 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c155
*+ bl_0_155 br_0_155 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c155
*+ bl_0_155 br_0_155 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c155
*+ bl_0_155 br_0_155 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c155
*+ bl_0_155 br_0_155 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c155
*+ bl_0_155 br_0_155 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c155
*+ bl_0_155 br_0_155 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c155
*+ bl_0_155 br_0_155 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c155
*+ bl_0_155 br_0_155 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c155
*+ bl_0_155 br_0_155 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c155
*+ bl_0_155 br_0_155 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c155
*+ bl_0_155 br_0_155 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c155
*+ bl_0_155 br_0_155 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c155
*+ bl_0_155 br_0_155 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c155
*+ bl_0_155 br_0_155 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c155
*+ bl_0_155 br_0_155 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c155
*+ bl_0_155 br_0_155 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c155
*+ bl_0_155 br_0_155 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c155
*+ bl_0_155 br_0_155 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c155
*+ bl_0_155 br_0_155 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c155
*+ bl_0_155 br_0_155 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c155
*+ bl_0_155 br_0_155 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c155
*+ bl_0_155 br_0_155 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c155
*+ bl_0_155 br_0_155 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c155
*+ bl_0_155 br_0_155 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c155
*+ bl_0_155 br_0_155 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c155
*+ bl_0_155 br_0_155 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c155
*+ bl_0_155 br_0_155 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c155
*+ bl_0_155 br_0_155 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c155
*+ bl_0_155 br_0_155 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c155
*+ bl_0_155 br_0_155 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c155
*+ bl_0_155 br_0_155 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c155
*+ bl_0_155 br_0_155 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c155
*+ bl_0_155 br_0_155 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c155
*+ bl_0_155 br_0_155 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c155
*+ bl_0_155 br_0_155 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c155
*+ bl_0_155 br_0_155 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c155
*+ bl_0_155 br_0_155 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c155
*+ bl_0_155 br_0_155 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c155
*+ bl_0_155 br_0_155 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c155
*+ bl_0_155 br_0_155 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c155
*+ bl_0_155 br_0_155 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c155
*+ bl_0_155 br_0_155 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c155
*+ bl_0_155 br_0_155 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c155
*+ bl_0_155 br_0_155 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c155
*+ bl_0_155 br_0_155 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c155
*+ bl_0_155 br_0_155 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c155
*+ bl_0_155 br_0_155 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c155
*+ bl_0_155 br_0_155 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c155
*+ bl_0_155 br_0_155 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c155
*+ bl_0_155 br_0_155 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c155
*+ bl_0_155 br_0_155 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c155
*+ bl_0_155 br_0_155 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c155
*+ bl_0_155 br_0_155 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c155
*+ bl_0_155 br_0_155 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c155
*+ bl_0_155 br_0_155 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c155
*+ bl_0_155 br_0_155 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c155
*+ bl_0_155 br_0_155 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c155
*+ bl_0_155 br_0_155 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c155
*+ bl_0_155 br_0_155 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c155
*+ bl_0_155 br_0_155 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c155
*+ bl_0_155 br_0_155 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c155
*+ bl_0_155 br_0_155 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c155
*+ bl_0_155 br_0_155 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c155
*+ bl_0_155 br_0_155 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c155
*+ bl_0_155 br_0_155 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c155
*+ bl_0_155 br_0_155 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c155
*+ bl_0_155 br_0_155 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c155
*+ bl_0_155 br_0_155 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c155
*+ bl_0_155 br_0_155 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c155
*+ bl_0_155 br_0_155 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c155
*+ bl_0_155 br_0_155 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c155
*+ bl_0_155 br_0_155 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c155
*+ bl_0_155 br_0_155 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c155
*+ bl_0_155 br_0_155 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c155
*+ bl_0_155 br_0_155 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c155
*+ bl_0_155 br_0_155 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c155
*+ bl_0_155 br_0_155 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c155
*+ bl_0_155 br_0_155 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c155
*+ bl_0_155 br_0_155 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c155
*+ bl_0_155 br_0_155 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c155
*+ bl_0_155 br_0_155 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c155
*+ bl_0_155 br_0_155 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c155
*+ bl_0_155 br_0_155 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c155
*+ bl_0_155 br_0_155 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c155
*+ bl_0_155 br_0_155 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c155
*+ bl_0_155 br_0_155 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c155
*+ bl_0_155 br_0_155 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c155
*+ bl_0_155 br_0_155 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c155
*+ bl_0_155 br_0_155 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c155
*+ bl_0_155 br_0_155 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c155
*+ bl_0_155 br_0_155 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c155
*+ bl_0_155 br_0_155 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c155
*+ bl_0_155 br_0_155 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c155
*+ bl_0_155 br_0_155 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c155
*+ bl_0_155 br_0_155 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c155
+ bl_0_155 br_0_155 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c156
+ bl_0_156 br_0_156 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c156
*+ bl_0_156 br_0_156 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c156
*+ bl_0_156 br_0_156 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c156
*+ bl_0_156 br_0_156 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c156
*+ bl_0_156 br_0_156 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c156
*+ bl_0_156 br_0_156 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c156
*+ bl_0_156 br_0_156 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c156
*+ bl_0_156 br_0_156 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c156
*+ bl_0_156 br_0_156 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c156
*+ bl_0_156 br_0_156 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c156
*+ bl_0_156 br_0_156 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c156
*+ bl_0_156 br_0_156 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c156
*+ bl_0_156 br_0_156 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c156
*+ bl_0_156 br_0_156 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c156
*+ bl_0_156 br_0_156 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c156
*+ bl_0_156 br_0_156 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c156
*+ bl_0_156 br_0_156 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c156
*+ bl_0_156 br_0_156 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c156
*+ bl_0_156 br_0_156 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c156
*+ bl_0_156 br_0_156 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c156
*+ bl_0_156 br_0_156 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c156
*+ bl_0_156 br_0_156 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c156
*+ bl_0_156 br_0_156 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c156
*+ bl_0_156 br_0_156 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c156
*+ bl_0_156 br_0_156 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c156
*+ bl_0_156 br_0_156 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c156
*+ bl_0_156 br_0_156 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c156
*+ bl_0_156 br_0_156 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c156
*+ bl_0_156 br_0_156 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c156
*+ bl_0_156 br_0_156 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c156
*+ bl_0_156 br_0_156 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c156
*+ bl_0_156 br_0_156 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c156
*+ bl_0_156 br_0_156 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c156
*+ bl_0_156 br_0_156 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c156
*+ bl_0_156 br_0_156 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c156
*+ bl_0_156 br_0_156 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c156
*+ bl_0_156 br_0_156 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c156
*+ bl_0_156 br_0_156 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c156
*+ bl_0_156 br_0_156 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c156
*+ bl_0_156 br_0_156 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c156
*+ bl_0_156 br_0_156 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c156
*+ bl_0_156 br_0_156 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c156
*+ bl_0_156 br_0_156 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c156
*+ bl_0_156 br_0_156 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c156
*+ bl_0_156 br_0_156 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c156
*+ bl_0_156 br_0_156 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c156
*+ bl_0_156 br_0_156 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c156
*+ bl_0_156 br_0_156 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c156
*+ bl_0_156 br_0_156 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c156
*+ bl_0_156 br_0_156 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c156
*+ bl_0_156 br_0_156 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c156
*+ bl_0_156 br_0_156 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c156
*+ bl_0_156 br_0_156 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c156
*+ bl_0_156 br_0_156 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c156
*+ bl_0_156 br_0_156 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c156
*+ bl_0_156 br_0_156 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c156
*+ bl_0_156 br_0_156 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c156
*+ bl_0_156 br_0_156 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c156
*+ bl_0_156 br_0_156 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c156
*+ bl_0_156 br_0_156 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c156
*+ bl_0_156 br_0_156 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c156
*+ bl_0_156 br_0_156 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c156
*+ bl_0_156 br_0_156 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c156
*+ bl_0_156 br_0_156 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c156
*+ bl_0_156 br_0_156 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c156
*+ bl_0_156 br_0_156 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c156
*+ bl_0_156 br_0_156 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c156
*+ bl_0_156 br_0_156 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c156
*+ bl_0_156 br_0_156 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c156
*+ bl_0_156 br_0_156 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c156
*+ bl_0_156 br_0_156 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c156
*+ bl_0_156 br_0_156 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c156
*+ bl_0_156 br_0_156 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c156
*+ bl_0_156 br_0_156 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c156
*+ bl_0_156 br_0_156 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c156
*+ bl_0_156 br_0_156 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c156
*+ bl_0_156 br_0_156 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c156
*+ bl_0_156 br_0_156 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c156
*+ bl_0_156 br_0_156 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c156
*+ bl_0_156 br_0_156 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c156
*+ bl_0_156 br_0_156 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c156
*+ bl_0_156 br_0_156 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c156
*+ bl_0_156 br_0_156 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c156
*+ bl_0_156 br_0_156 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c156
*+ bl_0_156 br_0_156 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c156
*+ bl_0_156 br_0_156 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c156
*+ bl_0_156 br_0_156 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c156
*+ bl_0_156 br_0_156 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c156
*+ bl_0_156 br_0_156 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c156
*+ bl_0_156 br_0_156 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c156
*+ bl_0_156 br_0_156 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c156
*+ bl_0_156 br_0_156 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c156
*+ bl_0_156 br_0_156 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c156
*+ bl_0_156 br_0_156 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c156
*+ bl_0_156 br_0_156 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c156
*+ bl_0_156 br_0_156 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c156
*+ bl_0_156 br_0_156 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c156
*+ bl_0_156 br_0_156 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c156
*+ bl_0_156 br_0_156 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c156
*+ bl_0_156 br_0_156 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c156
*+ bl_0_156 br_0_156 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c156
*+ bl_0_156 br_0_156 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c156
*+ bl_0_156 br_0_156 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c156
*+ bl_0_156 br_0_156 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c156
*+ bl_0_156 br_0_156 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c156
*+ bl_0_156 br_0_156 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c156
*+ bl_0_156 br_0_156 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c156
*+ bl_0_156 br_0_156 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c156
*+ bl_0_156 br_0_156 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c156
*+ bl_0_156 br_0_156 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c156
*+ bl_0_156 br_0_156 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c156
*+ bl_0_156 br_0_156 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c156
*+ bl_0_156 br_0_156 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c156
*+ bl_0_156 br_0_156 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c156
*+ bl_0_156 br_0_156 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c156
*+ bl_0_156 br_0_156 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c156
*+ bl_0_156 br_0_156 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c156
*+ bl_0_156 br_0_156 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c156
*+ bl_0_156 br_0_156 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c156
*+ bl_0_156 br_0_156 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c156
*+ bl_0_156 br_0_156 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c156
*+ bl_0_156 br_0_156 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c156
*+ bl_0_156 br_0_156 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c156
*+ bl_0_156 br_0_156 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c156
*+ bl_0_156 br_0_156 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c156
*+ bl_0_156 br_0_156 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c156
*+ bl_0_156 br_0_156 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c156
+ bl_0_156 br_0_156 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c157
+ bl_0_157 br_0_157 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c157
*+ bl_0_157 br_0_157 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c157
*+ bl_0_157 br_0_157 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c157
*+ bl_0_157 br_0_157 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c157
*+ bl_0_157 br_0_157 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c157
*+ bl_0_157 br_0_157 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c157
*+ bl_0_157 br_0_157 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c157
*+ bl_0_157 br_0_157 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c157
*+ bl_0_157 br_0_157 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c157
*+ bl_0_157 br_0_157 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c157
*+ bl_0_157 br_0_157 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c157
*+ bl_0_157 br_0_157 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c157
*+ bl_0_157 br_0_157 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c157
*+ bl_0_157 br_0_157 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c157
*+ bl_0_157 br_0_157 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c157
*+ bl_0_157 br_0_157 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c157
*+ bl_0_157 br_0_157 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c157
*+ bl_0_157 br_0_157 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c157
*+ bl_0_157 br_0_157 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c157
*+ bl_0_157 br_0_157 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c157
*+ bl_0_157 br_0_157 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c157
*+ bl_0_157 br_0_157 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c157
*+ bl_0_157 br_0_157 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c157
*+ bl_0_157 br_0_157 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c157
*+ bl_0_157 br_0_157 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c157
*+ bl_0_157 br_0_157 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c157
*+ bl_0_157 br_0_157 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c157
*+ bl_0_157 br_0_157 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c157
*+ bl_0_157 br_0_157 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c157
*+ bl_0_157 br_0_157 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c157
*+ bl_0_157 br_0_157 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c157
*+ bl_0_157 br_0_157 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c157
*+ bl_0_157 br_0_157 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c157
*+ bl_0_157 br_0_157 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c157
*+ bl_0_157 br_0_157 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c157
*+ bl_0_157 br_0_157 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c157
*+ bl_0_157 br_0_157 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c157
*+ bl_0_157 br_0_157 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c157
*+ bl_0_157 br_0_157 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c157
*+ bl_0_157 br_0_157 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c157
*+ bl_0_157 br_0_157 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c157
*+ bl_0_157 br_0_157 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c157
*+ bl_0_157 br_0_157 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c157
*+ bl_0_157 br_0_157 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c157
*+ bl_0_157 br_0_157 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c157
*+ bl_0_157 br_0_157 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c157
*+ bl_0_157 br_0_157 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c157
*+ bl_0_157 br_0_157 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c157
*+ bl_0_157 br_0_157 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c157
*+ bl_0_157 br_0_157 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c157
*+ bl_0_157 br_0_157 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c157
*+ bl_0_157 br_0_157 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c157
*+ bl_0_157 br_0_157 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c157
*+ bl_0_157 br_0_157 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c157
*+ bl_0_157 br_0_157 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c157
*+ bl_0_157 br_0_157 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c157
*+ bl_0_157 br_0_157 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c157
*+ bl_0_157 br_0_157 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c157
*+ bl_0_157 br_0_157 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c157
*+ bl_0_157 br_0_157 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c157
*+ bl_0_157 br_0_157 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c157
*+ bl_0_157 br_0_157 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c157
*+ bl_0_157 br_0_157 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c157
*+ bl_0_157 br_0_157 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c157
*+ bl_0_157 br_0_157 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c157
*+ bl_0_157 br_0_157 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c157
*+ bl_0_157 br_0_157 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c157
*+ bl_0_157 br_0_157 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c157
*+ bl_0_157 br_0_157 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c157
*+ bl_0_157 br_0_157 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c157
*+ bl_0_157 br_0_157 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c157
*+ bl_0_157 br_0_157 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c157
*+ bl_0_157 br_0_157 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c157
*+ bl_0_157 br_0_157 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c157
*+ bl_0_157 br_0_157 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c157
*+ bl_0_157 br_0_157 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c157
*+ bl_0_157 br_0_157 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c157
*+ bl_0_157 br_0_157 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c157
*+ bl_0_157 br_0_157 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c157
*+ bl_0_157 br_0_157 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c157
*+ bl_0_157 br_0_157 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c157
*+ bl_0_157 br_0_157 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c157
*+ bl_0_157 br_0_157 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c157
*+ bl_0_157 br_0_157 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c157
*+ bl_0_157 br_0_157 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c157
*+ bl_0_157 br_0_157 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c157
*+ bl_0_157 br_0_157 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c157
*+ bl_0_157 br_0_157 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c157
*+ bl_0_157 br_0_157 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c157
*+ bl_0_157 br_0_157 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c157
*+ bl_0_157 br_0_157 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c157
*+ bl_0_157 br_0_157 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c157
*+ bl_0_157 br_0_157 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c157
*+ bl_0_157 br_0_157 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c157
*+ bl_0_157 br_0_157 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c157
*+ bl_0_157 br_0_157 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c157
*+ bl_0_157 br_0_157 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c157
*+ bl_0_157 br_0_157 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c157
*+ bl_0_157 br_0_157 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c157
*+ bl_0_157 br_0_157 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c157
*+ bl_0_157 br_0_157 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c157
*+ bl_0_157 br_0_157 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c157
*+ bl_0_157 br_0_157 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c157
*+ bl_0_157 br_0_157 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c157
*+ bl_0_157 br_0_157 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c157
*+ bl_0_157 br_0_157 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c157
*+ bl_0_157 br_0_157 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c157
*+ bl_0_157 br_0_157 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c157
*+ bl_0_157 br_0_157 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c157
*+ bl_0_157 br_0_157 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c157
*+ bl_0_157 br_0_157 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c157
*+ bl_0_157 br_0_157 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c157
*+ bl_0_157 br_0_157 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c157
*+ bl_0_157 br_0_157 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c157
*+ bl_0_157 br_0_157 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c157
*+ bl_0_157 br_0_157 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c157
*+ bl_0_157 br_0_157 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c157
*+ bl_0_157 br_0_157 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c157
*+ bl_0_157 br_0_157 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c157
*+ bl_0_157 br_0_157 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c157
*+ bl_0_157 br_0_157 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c157
*+ bl_0_157 br_0_157 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c157
*+ bl_0_157 br_0_157 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c157
*+ bl_0_157 br_0_157 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c157
*+ bl_0_157 br_0_157 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c157
*+ bl_0_157 br_0_157 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c157
*+ bl_0_157 br_0_157 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c157
+ bl_0_157 br_0_157 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c158
+ bl_0_158 br_0_158 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c158
*+ bl_0_158 br_0_158 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c158
*+ bl_0_158 br_0_158 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c158
*+ bl_0_158 br_0_158 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c158
*+ bl_0_158 br_0_158 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c158
*+ bl_0_158 br_0_158 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c158
*+ bl_0_158 br_0_158 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c158
*+ bl_0_158 br_0_158 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c158
*+ bl_0_158 br_0_158 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c158
*+ bl_0_158 br_0_158 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c158
*+ bl_0_158 br_0_158 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c158
*+ bl_0_158 br_0_158 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c158
*+ bl_0_158 br_0_158 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c158
*+ bl_0_158 br_0_158 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c158
*+ bl_0_158 br_0_158 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c158
*+ bl_0_158 br_0_158 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c158
*+ bl_0_158 br_0_158 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c158
*+ bl_0_158 br_0_158 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c158
*+ bl_0_158 br_0_158 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c158
*+ bl_0_158 br_0_158 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c158
*+ bl_0_158 br_0_158 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c158
*+ bl_0_158 br_0_158 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c158
*+ bl_0_158 br_0_158 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c158
*+ bl_0_158 br_0_158 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c158
*+ bl_0_158 br_0_158 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c158
*+ bl_0_158 br_0_158 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c158
*+ bl_0_158 br_0_158 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c158
*+ bl_0_158 br_0_158 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c158
*+ bl_0_158 br_0_158 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c158
*+ bl_0_158 br_0_158 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c158
*+ bl_0_158 br_0_158 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c158
*+ bl_0_158 br_0_158 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c158
*+ bl_0_158 br_0_158 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c158
*+ bl_0_158 br_0_158 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c158
*+ bl_0_158 br_0_158 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c158
*+ bl_0_158 br_0_158 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c158
*+ bl_0_158 br_0_158 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c158
*+ bl_0_158 br_0_158 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c158
*+ bl_0_158 br_0_158 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c158
*+ bl_0_158 br_0_158 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c158
*+ bl_0_158 br_0_158 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c158
*+ bl_0_158 br_0_158 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c158
*+ bl_0_158 br_0_158 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c158
*+ bl_0_158 br_0_158 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c158
*+ bl_0_158 br_0_158 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c158
*+ bl_0_158 br_0_158 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c158
*+ bl_0_158 br_0_158 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c158
*+ bl_0_158 br_0_158 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c158
*+ bl_0_158 br_0_158 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c158
*+ bl_0_158 br_0_158 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c158
*+ bl_0_158 br_0_158 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c158
*+ bl_0_158 br_0_158 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c158
*+ bl_0_158 br_0_158 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c158
*+ bl_0_158 br_0_158 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c158
*+ bl_0_158 br_0_158 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c158
*+ bl_0_158 br_0_158 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c158
*+ bl_0_158 br_0_158 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c158
*+ bl_0_158 br_0_158 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c158
*+ bl_0_158 br_0_158 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c158
*+ bl_0_158 br_0_158 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c158
*+ bl_0_158 br_0_158 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c158
*+ bl_0_158 br_0_158 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c158
*+ bl_0_158 br_0_158 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c158
*+ bl_0_158 br_0_158 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c158
*+ bl_0_158 br_0_158 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c158
*+ bl_0_158 br_0_158 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c158
*+ bl_0_158 br_0_158 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c158
*+ bl_0_158 br_0_158 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c158
*+ bl_0_158 br_0_158 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c158
*+ bl_0_158 br_0_158 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c158
*+ bl_0_158 br_0_158 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c158
*+ bl_0_158 br_0_158 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c158
*+ bl_0_158 br_0_158 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c158
*+ bl_0_158 br_0_158 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c158
*+ bl_0_158 br_0_158 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c158
*+ bl_0_158 br_0_158 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c158
*+ bl_0_158 br_0_158 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c158
*+ bl_0_158 br_0_158 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c158
*+ bl_0_158 br_0_158 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c158
*+ bl_0_158 br_0_158 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c158
*+ bl_0_158 br_0_158 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c158
*+ bl_0_158 br_0_158 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c158
*+ bl_0_158 br_0_158 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c158
*+ bl_0_158 br_0_158 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c158
*+ bl_0_158 br_0_158 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c158
*+ bl_0_158 br_0_158 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c158
*+ bl_0_158 br_0_158 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c158
*+ bl_0_158 br_0_158 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c158
*+ bl_0_158 br_0_158 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c158
*+ bl_0_158 br_0_158 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c158
*+ bl_0_158 br_0_158 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c158
*+ bl_0_158 br_0_158 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c158
*+ bl_0_158 br_0_158 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c158
*+ bl_0_158 br_0_158 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c158
*+ bl_0_158 br_0_158 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c158
*+ bl_0_158 br_0_158 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c158
*+ bl_0_158 br_0_158 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c158
*+ bl_0_158 br_0_158 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c158
*+ bl_0_158 br_0_158 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c158
*+ bl_0_158 br_0_158 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c158
*+ bl_0_158 br_0_158 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c158
*+ bl_0_158 br_0_158 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c158
*+ bl_0_158 br_0_158 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c158
*+ bl_0_158 br_0_158 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c158
*+ bl_0_158 br_0_158 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c158
*+ bl_0_158 br_0_158 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c158
*+ bl_0_158 br_0_158 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c158
*+ bl_0_158 br_0_158 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c158
*+ bl_0_158 br_0_158 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c158
*+ bl_0_158 br_0_158 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c158
*+ bl_0_158 br_0_158 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c158
*+ bl_0_158 br_0_158 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c158
*+ bl_0_158 br_0_158 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c158
*+ bl_0_158 br_0_158 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c158
*+ bl_0_158 br_0_158 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c158
*+ bl_0_158 br_0_158 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c158
*+ bl_0_158 br_0_158 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c158
*+ bl_0_158 br_0_158 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c158
*+ bl_0_158 br_0_158 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c158
*+ bl_0_158 br_0_158 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c158
*+ bl_0_158 br_0_158 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c158
*+ bl_0_158 br_0_158 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c158
*+ bl_0_158 br_0_158 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c158
*+ bl_0_158 br_0_158 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c158
*+ bl_0_158 br_0_158 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c158
*+ bl_0_158 br_0_158 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c158
*+ bl_0_158 br_0_158 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c158
+ bl_0_158 br_0_158 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c159
+ bl_0_159 br_0_159 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c159
*+ bl_0_159 br_0_159 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c159
*+ bl_0_159 br_0_159 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c159
*+ bl_0_159 br_0_159 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c159
*+ bl_0_159 br_0_159 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c159
*+ bl_0_159 br_0_159 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c159
*+ bl_0_159 br_0_159 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c159
*+ bl_0_159 br_0_159 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c159
*+ bl_0_159 br_0_159 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c159
*+ bl_0_159 br_0_159 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c159
*+ bl_0_159 br_0_159 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c159
*+ bl_0_159 br_0_159 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c159
*+ bl_0_159 br_0_159 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c159
*+ bl_0_159 br_0_159 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c159
*+ bl_0_159 br_0_159 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c159
*+ bl_0_159 br_0_159 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c159
*+ bl_0_159 br_0_159 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c159
*+ bl_0_159 br_0_159 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c159
*+ bl_0_159 br_0_159 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c159
*+ bl_0_159 br_0_159 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c159
*+ bl_0_159 br_0_159 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c159
*+ bl_0_159 br_0_159 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c159
*+ bl_0_159 br_0_159 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c159
*+ bl_0_159 br_0_159 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c159
*+ bl_0_159 br_0_159 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c159
*+ bl_0_159 br_0_159 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c159
*+ bl_0_159 br_0_159 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c159
*+ bl_0_159 br_0_159 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c159
*+ bl_0_159 br_0_159 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c159
*+ bl_0_159 br_0_159 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c159
*+ bl_0_159 br_0_159 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c159
*+ bl_0_159 br_0_159 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c159
*+ bl_0_159 br_0_159 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c159
*+ bl_0_159 br_0_159 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c159
*+ bl_0_159 br_0_159 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c159
*+ bl_0_159 br_0_159 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c159
*+ bl_0_159 br_0_159 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c159
*+ bl_0_159 br_0_159 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c159
*+ bl_0_159 br_0_159 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c159
*+ bl_0_159 br_0_159 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c159
*+ bl_0_159 br_0_159 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c159
*+ bl_0_159 br_0_159 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c159
*+ bl_0_159 br_0_159 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c159
*+ bl_0_159 br_0_159 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c159
*+ bl_0_159 br_0_159 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c159
*+ bl_0_159 br_0_159 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c159
*+ bl_0_159 br_0_159 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c159
*+ bl_0_159 br_0_159 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c159
*+ bl_0_159 br_0_159 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c159
*+ bl_0_159 br_0_159 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c159
*+ bl_0_159 br_0_159 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c159
*+ bl_0_159 br_0_159 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c159
*+ bl_0_159 br_0_159 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c159
*+ bl_0_159 br_0_159 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c159
*+ bl_0_159 br_0_159 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c159
*+ bl_0_159 br_0_159 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c159
*+ bl_0_159 br_0_159 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c159
*+ bl_0_159 br_0_159 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c159
*+ bl_0_159 br_0_159 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c159
*+ bl_0_159 br_0_159 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c159
*+ bl_0_159 br_0_159 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c159
*+ bl_0_159 br_0_159 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c159
*+ bl_0_159 br_0_159 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c159
*+ bl_0_159 br_0_159 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c159
*+ bl_0_159 br_0_159 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c159
*+ bl_0_159 br_0_159 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c159
*+ bl_0_159 br_0_159 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c159
*+ bl_0_159 br_0_159 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c159
*+ bl_0_159 br_0_159 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c159
*+ bl_0_159 br_0_159 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c159
*+ bl_0_159 br_0_159 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c159
*+ bl_0_159 br_0_159 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c159
*+ bl_0_159 br_0_159 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c159
*+ bl_0_159 br_0_159 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c159
*+ bl_0_159 br_0_159 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c159
*+ bl_0_159 br_0_159 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c159
*+ bl_0_159 br_0_159 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c159
*+ bl_0_159 br_0_159 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c159
*+ bl_0_159 br_0_159 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c159
*+ bl_0_159 br_0_159 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c159
*+ bl_0_159 br_0_159 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c159
*+ bl_0_159 br_0_159 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c159
*+ bl_0_159 br_0_159 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c159
*+ bl_0_159 br_0_159 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c159
*+ bl_0_159 br_0_159 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c159
*+ bl_0_159 br_0_159 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c159
*+ bl_0_159 br_0_159 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c159
*+ bl_0_159 br_0_159 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c159
*+ bl_0_159 br_0_159 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c159
*+ bl_0_159 br_0_159 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c159
*+ bl_0_159 br_0_159 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c159
*+ bl_0_159 br_0_159 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c159
*+ bl_0_159 br_0_159 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c159
*+ bl_0_159 br_0_159 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c159
*+ bl_0_159 br_0_159 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c159
*+ bl_0_159 br_0_159 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c159
*+ bl_0_159 br_0_159 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c159
*+ bl_0_159 br_0_159 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c159
*+ bl_0_159 br_0_159 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c159
*+ bl_0_159 br_0_159 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c159
*+ bl_0_159 br_0_159 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c159
*+ bl_0_159 br_0_159 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c159
*+ bl_0_159 br_0_159 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c159
*+ bl_0_159 br_0_159 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c159
*+ bl_0_159 br_0_159 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c159
*+ bl_0_159 br_0_159 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c159
*+ bl_0_159 br_0_159 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c159
*+ bl_0_159 br_0_159 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c159
*+ bl_0_159 br_0_159 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c159
*+ bl_0_159 br_0_159 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c159
*+ bl_0_159 br_0_159 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c159
*+ bl_0_159 br_0_159 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c159
*+ bl_0_159 br_0_159 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c159
*+ bl_0_159 br_0_159 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c159
*+ bl_0_159 br_0_159 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c159
*+ bl_0_159 br_0_159 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c159
*+ bl_0_159 br_0_159 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c159
*+ bl_0_159 br_0_159 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c159
*+ bl_0_159 br_0_159 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c159
*+ bl_0_159 br_0_159 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c159
*+ bl_0_159 br_0_159 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c159
*+ bl_0_159 br_0_159 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c159
*+ bl_0_159 br_0_159 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c159
*+ bl_0_159 br_0_159 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c159
*+ bl_0_159 br_0_159 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c159
*+ bl_0_159 br_0_159 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c159
*+ bl_0_159 br_0_159 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c159
+ bl_0_159 br_0_159 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c160
+ bl_0_160 br_0_160 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c160
*+ bl_0_160 br_0_160 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c160
*+ bl_0_160 br_0_160 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c160
*+ bl_0_160 br_0_160 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c160
*+ bl_0_160 br_0_160 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c160
*+ bl_0_160 br_0_160 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c160
*+ bl_0_160 br_0_160 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c160
*+ bl_0_160 br_0_160 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c160
*+ bl_0_160 br_0_160 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c160
*+ bl_0_160 br_0_160 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c160
*+ bl_0_160 br_0_160 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c160
*+ bl_0_160 br_0_160 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c160
*+ bl_0_160 br_0_160 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c160
*+ bl_0_160 br_0_160 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c160
*+ bl_0_160 br_0_160 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c160
*+ bl_0_160 br_0_160 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c160
*+ bl_0_160 br_0_160 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c160
*+ bl_0_160 br_0_160 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c160
*+ bl_0_160 br_0_160 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c160
*+ bl_0_160 br_0_160 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c160
*+ bl_0_160 br_0_160 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c160
*+ bl_0_160 br_0_160 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c160
*+ bl_0_160 br_0_160 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c160
*+ bl_0_160 br_0_160 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c160
*+ bl_0_160 br_0_160 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c160
*+ bl_0_160 br_0_160 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c160
*+ bl_0_160 br_0_160 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c160
*+ bl_0_160 br_0_160 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c160
*+ bl_0_160 br_0_160 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c160
*+ bl_0_160 br_0_160 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c160
*+ bl_0_160 br_0_160 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c160
*+ bl_0_160 br_0_160 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c160
*+ bl_0_160 br_0_160 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c160
*+ bl_0_160 br_0_160 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c160
*+ bl_0_160 br_0_160 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c160
*+ bl_0_160 br_0_160 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c160
*+ bl_0_160 br_0_160 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c160
*+ bl_0_160 br_0_160 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c160
*+ bl_0_160 br_0_160 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c160
*+ bl_0_160 br_0_160 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c160
*+ bl_0_160 br_0_160 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c160
*+ bl_0_160 br_0_160 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c160
*+ bl_0_160 br_0_160 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c160
*+ bl_0_160 br_0_160 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c160
*+ bl_0_160 br_0_160 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c160
*+ bl_0_160 br_0_160 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c160
*+ bl_0_160 br_0_160 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c160
*+ bl_0_160 br_0_160 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c160
*+ bl_0_160 br_0_160 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c160
*+ bl_0_160 br_0_160 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c160
*+ bl_0_160 br_0_160 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c160
*+ bl_0_160 br_0_160 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c160
*+ bl_0_160 br_0_160 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c160
*+ bl_0_160 br_0_160 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c160
*+ bl_0_160 br_0_160 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c160
*+ bl_0_160 br_0_160 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c160
*+ bl_0_160 br_0_160 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c160
*+ bl_0_160 br_0_160 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c160
*+ bl_0_160 br_0_160 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c160
*+ bl_0_160 br_0_160 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c160
*+ bl_0_160 br_0_160 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c160
*+ bl_0_160 br_0_160 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c160
*+ bl_0_160 br_0_160 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c160
*+ bl_0_160 br_0_160 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c160
*+ bl_0_160 br_0_160 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c160
*+ bl_0_160 br_0_160 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c160
*+ bl_0_160 br_0_160 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c160
*+ bl_0_160 br_0_160 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c160
*+ bl_0_160 br_0_160 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c160
*+ bl_0_160 br_0_160 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c160
*+ bl_0_160 br_0_160 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c160
*+ bl_0_160 br_0_160 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c160
*+ bl_0_160 br_0_160 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c160
*+ bl_0_160 br_0_160 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c160
*+ bl_0_160 br_0_160 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c160
*+ bl_0_160 br_0_160 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c160
*+ bl_0_160 br_0_160 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c160
*+ bl_0_160 br_0_160 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c160
*+ bl_0_160 br_0_160 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c160
*+ bl_0_160 br_0_160 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c160
*+ bl_0_160 br_0_160 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c160
*+ bl_0_160 br_0_160 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c160
*+ bl_0_160 br_0_160 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c160
*+ bl_0_160 br_0_160 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c160
*+ bl_0_160 br_0_160 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c160
*+ bl_0_160 br_0_160 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c160
*+ bl_0_160 br_0_160 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c160
*+ bl_0_160 br_0_160 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c160
*+ bl_0_160 br_0_160 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c160
*+ bl_0_160 br_0_160 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c160
*+ bl_0_160 br_0_160 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c160
*+ bl_0_160 br_0_160 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c160
*+ bl_0_160 br_0_160 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c160
*+ bl_0_160 br_0_160 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c160
*+ bl_0_160 br_0_160 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c160
*+ bl_0_160 br_0_160 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c160
*+ bl_0_160 br_0_160 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c160
*+ bl_0_160 br_0_160 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c160
*+ bl_0_160 br_0_160 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c160
*+ bl_0_160 br_0_160 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c160
*+ bl_0_160 br_0_160 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c160
*+ bl_0_160 br_0_160 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c160
*+ bl_0_160 br_0_160 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c160
*+ bl_0_160 br_0_160 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c160
*+ bl_0_160 br_0_160 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c160
*+ bl_0_160 br_0_160 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c160
*+ bl_0_160 br_0_160 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c160
*+ bl_0_160 br_0_160 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c160
*+ bl_0_160 br_0_160 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c160
*+ bl_0_160 br_0_160 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c160
*+ bl_0_160 br_0_160 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c160
*+ bl_0_160 br_0_160 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c160
*+ bl_0_160 br_0_160 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c160
*+ bl_0_160 br_0_160 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c160
*+ bl_0_160 br_0_160 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c160
*+ bl_0_160 br_0_160 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c160
*+ bl_0_160 br_0_160 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c160
*+ bl_0_160 br_0_160 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c160
*+ bl_0_160 br_0_160 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c160
*+ bl_0_160 br_0_160 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c160
*+ bl_0_160 br_0_160 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c160
*+ bl_0_160 br_0_160 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c160
*+ bl_0_160 br_0_160 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c160
*+ bl_0_160 br_0_160 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c160
*+ bl_0_160 br_0_160 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c160
*+ bl_0_160 br_0_160 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c160
*+ bl_0_160 br_0_160 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c160
+ bl_0_160 br_0_160 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c161
+ bl_0_161 br_0_161 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c161
*+ bl_0_161 br_0_161 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c161
*+ bl_0_161 br_0_161 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c161
*+ bl_0_161 br_0_161 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c161
*+ bl_0_161 br_0_161 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c161
*+ bl_0_161 br_0_161 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c161
*+ bl_0_161 br_0_161 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c161
*+ bl_0_161 br_0_161 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c161
*+ bl_0_161 br_0_161 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c161
*+ bl_0_161 br_0_161 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c161
*+ bl_0_161 br_0_161 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c161
*+ bl_0_161 br_0_161 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c161
*+ bl_0_161 br_0_161 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c161
*+ bl_0_161 br_0_161 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c161
*+ bl_0_161 br_0_161 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c161
*+ bl_0_161 br_0_161 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c161
*+ bl_0_161 br_0_161 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c161
*+ bl_0_161 br_0_161 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c161
*+ bl_0_161 br_0_161 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c161
*+ bl_0_161 br_0_161 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c161
*+ bl_0_161 br_0_161 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c161
*+ bl_0_161 br_0_161 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c161
*+ bl_0_161 br_0_161 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c161
*+ bl_0_161 br_0_161 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c161
*+ bl_0_161 br_0_161 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c161
*+ bl_0_161 br_0_161 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c161
*+ bl_0_161 br_0_161 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c161
*+ bl_0_161 br_0_161 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c161
*+ bl_0_161 br_0_161 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c161
*+ bl_0_161 br_0_161 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c161
*+ bl_0_161 br_0_161 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c161
*+ bl_0_161 br_0_161 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c161
*+ bl_0_161 br_0_161 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c161
*+ bl_0_161 br_0_161 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c161
*+ bl_0_161 br_0_161 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c161
*+ bl_0_161 br_0_161 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c161
*+ bl_0_161 br_0_161 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c161
*+ bl_0_161 br_0_161 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c161
*+ bl_0_161 br_0_161 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c161
*+ bl_0_161 br_0_161 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c161
*+ bl_0_161 br_0_161 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c161
*+ bl_0_161 br_0_161 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c161
*+ bl_0_161 br_0_161 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c161
*+ bl_0_161 br_0_161 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c161
*+ bl_0_161 br_0_161 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c161
*+ bl_0_161 br_0_161 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c161
*+ bl_0_161 br_0_161 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c161
*+ bl_0_161 br_0_161 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c161
*+ bl_0_161 br_0_161 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c161
*+ bl_0_161 br_0_161 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c161
*+ bl_0_161 br_0_161 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c161
*+ bl_0_161 br_0_161 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c161
*+ bl_0_161 br_0_161 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c161
*+ bl_0_161 br_0_161 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c161
*+ bl_0_161 br_0_161 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c161
*+ bl_0_161 br_0_161 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c161
*+ bl_0_161 br_0_161 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c161
*+ bl_0_161 br_0_161 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c161
*+ bl_0_161 br_0_161 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c161
*+ bl_0_161 br_0_161 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c161
*+ bl_0_161 br_0_161 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c161
*+ bl_0_161 br_0_161 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c161
*+ bl_0_161 br_0_161 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c161
*+ bl_0_161 br_0_161 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c161
*+ bl_0_161 br_0_161 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c161
*+ bl_0_161 br_0_161 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c161
*+ bl_0_161 br_0_161 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c161
*+ bl_0_161 br_0_161 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c161
*+ bl_0_161 br_0_161 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c161
*+ bl_0_161 br_0_161 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c161
*+ bl_0_161 br_0_161 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c161
*+ bl_0_161 br_0_161 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c161
*+ bl_0_161 br_0_161 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c161
*+ bl_0_161 br_0_161 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c161
*+ bl_0_161 br_0_161 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c161
*+ bl_0_161 br_0_161 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c161
*+ bl_0_161 br_0_161 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c161
*+ bl_0_161 br_0_161 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c161
*+ bl_0_161 br_0_161 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c161
*+ bl_0_161 br_0_161 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c161
*+ bl_0_161 br_0_161 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c161
*+ bl_0_161 br_0_161 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c161
*+ bl_0_161 br_0_161 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c161
*+ bl_0_161 br_0_161 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c161
*+ bl_0_161 br_0_161 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c161
*+ bl_0_161 br_0_161 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c161
*+ bl_0_161 br_0_161 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c161
*+ bl_0_161 br_0_161 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c161
*+ bl_0_161 br_0_161 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c161
*+ bl_0_161 br_0_161 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c161
*+ bl_0_161 br_0_161 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c161
*+ bl_0_161 br_0_161 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c161
*+ bl_0_161 br_0_161 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c161
*+ bl_0_161 br_0_161 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c161
*+ bl_0_161 br_0_161 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c161
*+ bl_0_161 br_0_161 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c161
*+ bl_0_161 br_0_161 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c161
*+ bl_0_161 br_0_161 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c161
*+ bl_0_161 br_0_161 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c161
*+ bl_0_161 br_0_161 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c161
*+ bl_0_161 br_0_161 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c161
*+ bl_0_161 br_0_161 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c161
*+ bl_0_161 br_0_161 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c161
*+ bl_0_161 br_0_161 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c161
*+ bl_0_161 br_0_161 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c161
*+ bl_0_161 br_0_161 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c161
*+ bl_0_161 br_0_161 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c161
*+ bl_0_161 br_0_161 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c161
*+ bl_0_161 br_0_161 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c161
*+ bl_0_161 br_0_161 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c161
*+ bl_0_161 br_0_161 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c161
*+ bl_0_161 br_0_161 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c161
*+ bl_0_161 br_0_161 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c161
*+ bl_0_161 br_0_161 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c161
*+ bl_0_161 br_0_161 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c161
*+ bl_0_161 br_0_161 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c161
*+ bl_0_161 br_0_161 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c161
*+ bl_0_161 br_0_161 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c161
*+ bl_0_161 br_0_161 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c161
*+ bl_0_161 br_0_161 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c161
*+ bl_0_161 br_0_161 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c161
*+ bl_0_161 br_0_161 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c161
*+ bl_0_161 br_0_161 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c161
*+ bl_0_161 br_0_161 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c161
*+ bl_0_161 br_0_161 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c161
*+ bl_0_161 br_0_161 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c161
*+ bl_0_161 br_0_161 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c161
+ bl_0_161 br_0_161 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c162
+ bl_0_162 br_0_162 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c162
*+ bl_0_162 br_0_162 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c162
*+ bl_0_162 br_0_162 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c162
*+ bl_0_162 br_0_162 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c162
*+ bl_0_162 br_0_162 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c162
*+ bl_0_162 br_0_162 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c162
*+ bl_0_162 br_0_162 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c162
*+ bl_0_162 br_0_162 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c162
*+ bl_0_162 br_0_162 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c162
*+ bl_0_162 br_0_162 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c162
*+ bl_0_162 br_0_162 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c162
*+ bl_0_162 br_0_162 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c162
*+ bl_0_162 br_0_162 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c162
*+ bl_0_162 br_0_162 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c162
*+ bl_0_162 br_0_162 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c162
*+ bl_0_162 br_0_162 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c162
*+ bl_0_162 br_0_162 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c162
*+ bl_0_162 br_0_162 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c162
*+ bl_0_162 br_0_162 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c162
*+ bl_0_162 br_0_162 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c162
*+ bl_0_162 br_0_162 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c162
*+ bl_0_162 br_0_162 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c162
*+ bl_0_162 br_0_162 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c162
*+ bl_0_162 br_0_162 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c162
*+ bl_0_162 br_0_162 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c162
*+ bl_0_162 br_0_162 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c162
*+ bl_0_162 br_0_162 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c162
*+ bl_0_162 br_0_162 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c162
*+ bl_0_162 br_0_162 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c162
*+ bl_0_162 br_0_162 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c162
*+ bl_0_162 br_0_162 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c162
*+ bl_0_162 br_0_162 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c162
*+ bl_0_162 br_0_162 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c162
*+ bl_0_162 br_0_162 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c162
*+ bl_0_162 br_0_162 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c162
*+ bl_0_162 br_0_162 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c162
*+ bl_0_162 br_0_162 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c162
*+ bl_0_162 br_0_162 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c162
*+ bl_0_162 br_0_162 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c162
*+ bl_0_162 br_0_162 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c162
*+ bl_0_162 br_0_162 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c162
*+ bl_0_162 br_0_162 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c162
*+ bl_0_162 br_0_162 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c162
*+ bl_0_162 br_0_162 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c162
*+ bl_0_162 br_0_162 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c162
*+ bl_0_162 br_0_162 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c162
*+ bl_0_162 br_0_162 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c162
*+ bl_0_162 br_0_162 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c162
*+ bl_0_162 br_0_162 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c162
*+ bl_0_162 br_0_162 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c162
*+ bl_0_162 br_0_162 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c162
*+ bl_0_162 br_0_162 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c162
*+ bl_0_162 br_0_162 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c162
*+ bl_0_162 br_0_162 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c162
*+ bl_0_162 br_0_162 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c162
*+ bl_0_162 br_0_162 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c162
*+ bl_0_162 br_0_162 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c162
*+ bl_0_162 br_0_162 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c162
*+ bl_0_162 br_0_162 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c162
*+ bl_0_162 br_0_162 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c162
*+ bl_0_162 br_0_162 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c162
*+ bl_0_162 br_0_162 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c162
*+ bl_0_162 br_0_162 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c162
*+ bl_0_162 br_0_162 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c162
*+ bl_0_162 br_0_162 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c162
*+ bl_0_162 br_0_162 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c162
*+ bl_0_162 br_0_162 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c162
*+ bl_0_162 br_0_162 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c162
*+ bl_0_162 br_0_162 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c162
*+ bl_0_162 br_0_162 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c162
*+ bl_0_162 br_0_162 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c162
*+ bl_0_162 br_0_162 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c162
*+ bl_0_162 br_0_162 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c162
*+ bl_0_162 br_0_162 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c162
*+ bl_0_162 br_0_162 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c162
*+ bl_0_162 br_0_162 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c162
*+ bl_0_162 br_0_162 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c162
*+ bl_0_162 br_0_162 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c162
*+ bl_0_162 br_0_162 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c162
*+ bl_0_162 br_0_162 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c162
*+ bl_0_162 br_0_162 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c162
*+ bl_0_162 br_0_162 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c162
*+ bl_0_162 br_0_162 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c162
*+ bl_0_162 br_0_162 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c162
*+ bl_0_162 br_0_162 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c162
*+ bl_0_162 br_0_162 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c162
*+ bl_0_162 br_0_162 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c162
*+ bl_0_162 br_0_162 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c162
*+ bl_0_162 br_0_162 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c162
*+ bl_0_162 br_0_162 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c162
*+ bl_0_162 br_0_162 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c162
*+ bl_0_162 br_0_162 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c162
*+ bl_0_162 br_0_162 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c162
*+ bl_0_162 br_0_162 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c162
*+ bl_0_162 br_0_162 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c162
*+ bl_0_162 br_0_162 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c162
*+ bl_0_162 br_0_162 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c162
*+ bl_0_162 br_0_162 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c162
*+ bl_0_162 br_0_162 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c162
*+ bl_0_162 br_0_162 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c162
*+ bl_0_162 br_0_162 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c162
*+ bl_0_162 br_0_162 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c162
*+ bl_0_162 br_0_162 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c162
*+ bl_0_162 br_0_162 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c162
*+ bl_0_162 br_0_162 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c162
*+ bl_0_162 br_0_162 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c162
*+ bl_0_162 br_0_162 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c162
*+ bl_0_162 br_0_162 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c162
*+ bl_0_162 br_0_162 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c162
*+ bl_0_162 br_0_162 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c162
*+ bl_0_162 br_0_162 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c162
*+ bl_0_162 br_0_162 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c162
*+ bl_0_162 br_0_162 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c162
*+ bl_0_162 br_0_162 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c162
*+ bl_0_162 br_0_162 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c162
*+ bl_0_162 br_0_162 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c162
*+ bl_0_162 br_0_162 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c162
*+ bl_0_162 br_0_162 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c162
*+ bl_0_162 br_0_162 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c162
*+ bl_0_162 br_0_162 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c162
*+ bl_0_162 br_0_162 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c162
*+ bl_0_162 br_0_162 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c162
*+ bl_0_162 br_0_162 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c162
*+ bl_0_162 br_0_162 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c162
*+ bl_0_162 br_0_162 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c162
*+ bl_0_162 br_0_162 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c162
*+ bl_0_162 br_0_162 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c162
+ bl_0_162 br_0_162 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c163
+ bl_0_163 br_0_163 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c163
*+ bl_0_163 br_0_163 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c163
*+ bl_0_163 br_0_163 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c163
*+ bl_0_163 br_0_163 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c163
*+ bl_0_163 br_0_163 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c163
*+ bl_0_163 br_0_163 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c163
*+ bl_0_163 br_0_163 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c163
*+ bl_0_163 br_0_163 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c163
*+ bl_0_163 br_0_163 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c163
*+ bl_0_163 br_0_163 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c163
*+ bl_0_163 br_0_163 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c163
*+ bl_0_163 br_0_163 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c163
*+ bl_0_163 br_0_163 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c163
*+ bl_0_163 br_0_163 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c163
*+ bl_0_163 br_0_163 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c163
*+ bl_0_163 br_0_163 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c163
*+ bl_0_163 br_0_163 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c163
*+ bl_0_163 br_0_163 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c163
*+ bl_0_163 br_0_163 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c163
*+ bl_0_163 br_0_163 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c163
*+ bl_0_163 br_0_163 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c163
*+ bl_0_163 br_0_163 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c163
*+ bl_0_163 br_0_163 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c163
*+ bl_0_163 br_0_163 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c163
*+ bl_0_163 br_0_163 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c163
*+ bl_0_163 br_0_163 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c163
*+ bl_0_163 br_0_163 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c163
*+ bl_0_163 br_0_163 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c163
*+ bl_0_163 br_0_163 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c163
*+ bl_0_163 br_0_163 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c163
*+ bl_0_163 br_0_163 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c163
*+ bl_0_163 br_0_163 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c163
*+ bl_0_163 br_0_163 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c163
*+ bl_0_163 br_0_163 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c163
*+ bl_0_163 br_0_163 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c163
*+ bl_0_163 br_0_163 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c163
*+ bl_0_163 br_0_163 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c163
*+ bl_0_163 br_0_163 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c163
*+ bl_0_163 br_0_163 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c163
*+ bl_0_163 br_0_163 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c163
*+ bl_0_163 br_0_163 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c163
*+ bl_0_163 br_0_163 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c163
*+ bl_0_163 br_0_163 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c163
*+ bl_0_163 br_0_163 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c163
*+ bl_0_163 br_0_163 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c163
*+ bl_0_163 br_0_163 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c163
*+ bl_0_163 br_0_163 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c163
*+ bl_0_163 br_0_163 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c163
*+ bl_0_163 br_0_163 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c163
*+ bl_0_163 br_0_163 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c163
*+ bl_0_163 br_0_163 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c163
*+ bl_0_163 br_0_163 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c163
*+ bl_0_163 br_0_163 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c163
*+ bl_0_163 br_0_163 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c163
*+ bl_0_163 br_0_163 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c163
*+ bl_0_163 br_0_163 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c163
*+ bl_0_163 br_0_163 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c163
*+ bl_0_163 br_0_163 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c163
*+ bl_0_163 br_0_163 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c163
*+ bl_0_163 br_0_163 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c163
*+ bl_0_163 br_0_163 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c163
*+ bl_0_163 br_0_163 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c163
*+ bl_0_163 br_0_163 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c163
*+ bl_0_163 br_0_163 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c163
*+ bl_0_163 br_0_163 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c163
*+ bl_0_163 br_0_163 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c163
*+ bl_0_163 br_0_163 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c163
*+ bl_0_163 br_0_163 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c163
*+ bl_0_163 br_0_163 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c163
*+ bl_0_163 br_0_163 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c163
*+ bl_0_163 br_0_163 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c163
*+ bl_0_163 br_0_163 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c163
*+ bl_0_163 br_0_163 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c163
*+ bl_0_163 br_0_163 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c163
*+ bl_0_163 br_0_163 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c163
*+ bl_0_163 br_0_163 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c163
*+ bl_0_163 br_0_163 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c163
*+ bl_0_163 br_0_163 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c163
*+ bl_0_163 br_0_163 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c163
*+ bl_0_163 br_0_163 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c163
*+ bl_0_163 br_0_163 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c163
*+ bl_0_163 br_0_163 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c163
*+ bl_0_163 br_0_163 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c163
*+ bl_0_163 br_0_163 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c163
*+ bl_0_163 br_0_163 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c163
*+ bl_0_163 br_0_163 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c163
*+ bl_0_163 br_0_163 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c163
*+ bl_0_163 br_0_163 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c163
*+ bl_0_163 br_0_163 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c163
*+ bl_0_163 br_0_163 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c163
*+ bl_0_163 br_0_163 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c163
*+ bl_0_163 br_0_163 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c163
*+ bl_0_163 br_0_163 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c163
*+ bl_0_163 br_0_163 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c163
*+ bl_0_163 br_0_163 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c163
*+ bl_0_163 br_0_163 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c163
*+ bl_0_163 br_0_163 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c163
*+ bl_0_163 br_0_163 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c163
*+ bl_0_163 br_0_163 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c163
*+ bl_0_163 br_0_163 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c163
*+ bl_0_163 br_0_163 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c163
*+ bl_0_163 br_0_163 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c163
*+ bl_0_163 br_0_163 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c163
*+ bl_0_163 br_0_163 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c163
*+ bl_0_163 br_0_163 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c163
*+ bl_0_163 br_0_163 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c163
*+ bl_0_163 br_0_163 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c163
*+ bl_0_163 br_0_163 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c163
*+ bl_0_163 br_0_163 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c163
*+ bl_0_163 br_0_163 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c163
*+ bl_0_163 br_0_163 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c163
*+ bl_0_163 br_0_163 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c163
*+ bl_0_163 br_0_163 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c163
*+ bl_0_163 br_0_163 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c163
*+ bl_0_163 br_0_163 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c163
*+ bl_0_163 br_0_163 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c163
*+ bl_0_163 br_0_163 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c163
*+ bl_0_163 br_0_163 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c163
*+ bl_0_163 br_0_163 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c163
*+ bl_0_163 br_0_163 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c163
*+ bl_0_163 br_0_163 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c163
*+ bl_0_163 br_0_163 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c163
*+ bl_0_163 br_0_163 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c163
*+ bl_0_163 br_0_163 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c163
*+ bl_0_163 br_0_163 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c163
*+ bl_0_163 br_0_163 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c163
*+ bl_0_163 br_0_163 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c163
+ bl_0_163 br_0_163 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c164
+ bl_0_164 br_0_164 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c164
*+ bl_0_164 br_0_164 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c164
*+ bl_0_164 br_0_164 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c164
*+ bl_0_164 br_0_164 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c164
*+ bl_0_164 br_0_164 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c164
*+ bl_0_164 br_0_164 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c164
*+ bl_0_164 br_0_164 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c164
*+ bl_0_164 br_0_164 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c164
*+ bl_0_164 br_0_164 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c164
*+ bl_0_164 br_0_164 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c164
*+ bl_0_164 br_0_164 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c164
*+ bl_0_164 br_0_164 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c164
*+ bl_0_164 br_0_164 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c164
*+ bl_0_164 br_0_164 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c164
*+ bl_0_164 br_0_164 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c164
*+ bl_0_164 br_0_164 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c164
*+ bl_0_164 br_0_164 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c164
*+ bl_0_164 br_0_164 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c164
*+ bl_0_164 br_0_164 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c164
*+ bl_0_164 br_0_164 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c164
*+ bl_0_164 br_0_164 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c164
*+ bl_0_164 br_0_164 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c164
*+ bl_0_164 br_0_164 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c164
*+ bl_0_164 br_0_164 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c164
*+ bl_0_164 br_0_164 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c164
*+ bl_0_164 br_0_164 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c164
*+ bl_0_164 br_0_164 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c164
*+ bl_0_164 br_0_164 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c164
*+ bl_0_164 br_0_164 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c164
*+ bl_0_164 br_0_164 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c164
*+ bl_0_164 br_0_164 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c164
*+ bl_0_164 br_0_164 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c164
*+ bl_0_164 br_0_164 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c164
*+ bl_0_164 br_0_164 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c164
*+ bl_0_164 br_0_164 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c164
*+ bl_0_164 br_0_164 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c164
*+ bl_0_164 br_0_164 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c164
*+ bl_0_164 br_0_164 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c164
*+ bl_0_164 br_0_164 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c164
*+ bl_0_164 br_0_164 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c164
*+ bl_0_164 br_0_164 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c164
*+ bl_0_164 br_0_164 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c164
*+ bl_0_164 br_0_164 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c164
*+ bl_0_164 br_0_164 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c164
*+ bl_0_164 br_0_164 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c164
*+ bl_0_164 br_0_164 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c164
*+ bl_0_164 br_0_164 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c164
*+ bl_0_164 br_0_164 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c164
*+ bl_0_164 br_0_164 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c164
*+ bl_0_164 br_0_164 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c164
*+ bl_0_164 br_0_164 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c164
*+ bl_0_164 br_0_164 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c164
*+ bl_0_164 br_0_164 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c164
*+ bl_0_164 br_0_164 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c164
*+ bl_0_164 br_0_164 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c164
*+ bl_0_164 br_0_164 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c164
*+ bl_0_164 br_0_164 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c164
*+ bl_0_164 br_0_164 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c164
*+ bl_0_164 br_0_164 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c164
*+ bl_0_164 br_0_164 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c164
*+ bl_0_164 br_0_164 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c164
*+ bl_0_164 br_0_164 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c164
*+ bl_0_164 br_0_164 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c164
*+ bl_0_164 br_0_164 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c164
*+ bl_0_164 br_0_164 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c164
*+ bl_0_164 br_0_164 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c164
*+ bl_0_164 br_0_164 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c164
*+ bl_0_164 br_0_164 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c164
*+ bl_0_164 br_0_164 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c164
*+ bl_0_164 br_0_164 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c164
*+ bl_0_164 br_0_164 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c164
*+ bl_0_164 br_0_164 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c164
*+ bl_0_164 br_0_164 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c164
*+ bl_0_164 br_0_164 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c164
*+ bl_0_164 br_0_164 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c164
*+ bl_0_164 br_0_164 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c164
*+ bl_0_164 br_0_164 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c164
*+ bl_0_164 br_0_164 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c164
*+ bl_0_164 br_0_164 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c164
*+ bl_0_164 br_0_164 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c164
*+ bl_0_164 br_0_164 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c164
*+ bl_0_164 br_0_164 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c164
*+ bl_0_164 br_0_164 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c164
*+ bl_0_164 br_0_164 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c164
*+ bl_0_164 br_0_164 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c164
*+ bl_0_164 br_0_164 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c164
*+ bl_0_164 br_0_164 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c164
*+ bl_0_164 br_0_164 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c164
*+ bl_0_164 br_0_164 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c164
*+ bl_0_164 br_0_164 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c164
*+ bl_0_164 br_0_164 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c164
*+ bl_0_164 br_0_164 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c164
*+ bl_0_164 br_0_164 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c164
*+ bl_0_164 br_0_164 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c164
*+ bl_0_164 br_0_164 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c164
*+ bl_0_164 br_0_164 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c164
*+ bl_0_164 br_0_164 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c164
*+ bl_0_164 br_0_164 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c164
*+ bl_0_164 br_0_164 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c164
*+ bl_0_164 br_0_164 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c164
*+ bl_0_164 br_0_164 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c164
*+ bl_0_164 br_0_164 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c164
*+ bl_0_164 br_0_164 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c164
*+ bl_0_164 br_0_164 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c164
*+ bl_0_164 br_0_164 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c164
*+ bl_0_164 br_0_164 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c164
*+ bl_0_164 br_0_164 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c164
*+ bl_0_164 br_0_164 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c164
*+ bl_0_164 br_0_164 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c164
*+ bl_0_164 br_0_164 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c164
*+ bl_0_164 br_0_164 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c164
*+ bl_0_164 br_0_164 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c164
*+ bl_0_164 br_0_164 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c164
*+ bl_0_164 br_0_164 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c164
*+ bl_0_164 br_0_164 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c164
*+ bl_0_164 br_0_164 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c164
*+ bl_0_164 br_0_164 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c164
*+ bl_0_164 br_0_164 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c164
*+ bl_0_164 br_0_164 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c164
*+ bl_0_164 br_0_164 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c164
*+ bl_0_164 br_0_164 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c164
*+ bl_0_164 br_0_164 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c164
*+ bl_0_164 br_0_164 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c164
*+ bl_0_164 br_0_164 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c164
*+ bl_0_164 br_0_164 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c164
*+ bl_0_164 br_0_164 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c164
*+ bl_0_164 br_0_164 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c164
+ bl_0_164 br_0_164 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c165
+ bl_0_165 br_0_165 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c165
*+ bl_0_165 br_0_165 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c165
*+ bl_0_165 br_0_165 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c165
*+ bl_0_165 br_0_165 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c165
*+ bl_0_165 br_0_165 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c165
*+ bl_0_165 br_0_165 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c165
*+ bl_0_165 br_0_165 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c165
*+ bl_0_165 br_0_165 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c165
*+ bl_0_165 br_0_165 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c165
*+ bl_0_165 br_0_165 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c165
*+ bl_0_165 br_0_165 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c165
*+ bl_0_165 br_0_165 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c165
*+ bl_0_165 br_0_165 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c165
*+ bl_0_165 br_0_165 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c165
*+ bl_0_165 br_0_165 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c165
*+ bl_0_165 br_0_165 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c165
*+ bl_0_165 br_0_165 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c165
*+ bl_0_165 br_0_165 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c165
*+ bl_0_165 br_0_165 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c165
*+ bl_0_165 br_0_165 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c165
*+ bl_0_165 br_0_165 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c165
*+ bl_0_165 br_0_165 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c165
*+ bl_0_165 br_0_165 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c165
*+ bl_0_165 br_0_165 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c165
*+ bl_0_165 br_0_165 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c165
*+ bl_0_165 br_0_165 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c165
*+ bl_0_165 br_0_165 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c165
*+ bl_0_165 br_0_165 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c165
*+ bl_0_165 br_0_165 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c165
*+ bl_0_165 br_0_165 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c165
*+ bl_0_165 br_0_165 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c165
*+ bl_0_165 br_0_165 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c165
*+ bl_0_165 br_0_165 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c165
*+ bl_0_165 br_0_165 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c165
*+ bl_0_165 br_0_165 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c165
*+ bl_0_165 br_0_165 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c165
*+ bl_0_165 br_0_165 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c165
*+ bl_0_165 br_0_165 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c165
*+ bl_0_165 br_0_165 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c165
*+ bl_0_165 br_0_165 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c165
*+ bl_0_165 br_0_165 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c165
*+ bl_0_165 br_0_165 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c165
*+ bl_0_165 br_0_165 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c165
*+ bl_0_165 br_0_165 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c165
*+ bl_0_165 br_0_165 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c165
*+ bl_0_165 br_0_165 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c165
*+ bl_0_165 br_0_165 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c165
*+ bl_0_165 br_0_165 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c165
*+ bl_0_165 br_0_165 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c165
*+ bl_0_165 br_0_165 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c165
*+ bl_0_165 br_0_165 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c165
*+ bl_0_165 br_0_165 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c165
*+ bl_0_165 br_0_165 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c165
*+ bl_0_165 br_0_165 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c165
*+ bl_0_165 br_0_165 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c165
*+ bl_0_165 br_0_165 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c165
*+ bl_0_165 br_0_165 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c165
*+ bl_0_165 br_0_165 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c165
*+ bl_0_165 br_0_165 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c165
*+ bl_0_165 br_0_165 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c165
*+ bl_0_165 br_0_165 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c165
*+ bl_0_165 br_0_165 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c165
*+ bl_0_165 br_0_165 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c165
*+ bl_0_165 br_0_165 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c165
*+ bl_0_165 br_0_165 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c165
*+ bl_0_165 br_0_165 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c165
*+ bl_0_165 br_0_165 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c165
*+ bl_0_165 br_0_165 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c165
*+ bl_0_165 br_0_165 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c165
*+ bl_0_165 br_0_165 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c165
*+ bl_0_165 br_0_165 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c165
*+ bl_0_165 br_0_165 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c165
*+ bl_0_165 br_0_165 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c165
*+ bl_0_165 br_0_165 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c165
*+ bl_0_165 br_0_165 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c165
*+ bl_0_165 br_0_165 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c165
*+ bl_0_165 br_0_165 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c165
*+ bl_0_165 br_0_165 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c165
*+ bl_0_165 br_0_165 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c165
*+ bl_0_165 br_0_165 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c165
*+ bl_0_165 br_0_165 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c165
*+ bl_0_165 br_0_165 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c165
*+ bl_0_165 br_0_165 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c165
*+ bl_0_165 br_0_165 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c165
*+ bl_0_165 br_0_165 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c165
*+ bl_0_165 br_0_165 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c165
*+ bl_0_165 br_0_165 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c165
*+ bl_0_165 br_0_165 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c165
*+ bl_0_165 br_0_165 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c165
*+ bl_0_165 br_0_165 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c165
*+ bl_0_165 br_0_165 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c165
*+ bl_0_165 br_0_165 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c165
*+ bl_0_165 br_0_165 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c165
*+ bl_0_165 br_0_165 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c165
*+ bl_0_165 br_0_165 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c165
*+ bl_0_165 br_0_165 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c165
*+ bl_0_165 br_0_165 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c165
*+ bl_0_165 br_0_165 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c165
*+ bl_0_165 br_0_165 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c165
*+ bl_0_165 br_0_165 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c165
*+ bl_0_165 br_0_165 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c165
*+ bl_0_165 br_0_165 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c165
*+ bl_0_165 br_0_165 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c165
*+ bl_0_165 br_0_165 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c165
*+ bl_0_165 br_0_165 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c165
*+ bl_0_165 br_0_165 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c165
*+ bl_0_165 br_0_165 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c165
*+ bl_0_165 br_0_165 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c165
*+ bl_0_165 br_0_165 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c165
*+ bl_0_165 br_0_165 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c165
*+ bl_0_165 br_0_165 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c165
*+ bl_0_165 br_0_165 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c165
*+ bl_0_165 br_0_165 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c165
*+ bl_0_165 br_0_165 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c165
*+ bl_0_165 br_0_165 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c165
*+ bl_0_165 br_0_165 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c165
*+ bl_0_165 br_0_165 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c165
*+ bl_0_165 br_0_165 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c165
*+ bl_0_165 br_0_165 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c165
*+ bl_0_165 br_0_165 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c165
*+ bl_0_165 br_0_165 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c165
*+ bl_0_165 br_0_165 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c165
*+ bl_0_165 br_0_165 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c165
*+ bl_0_165 br_0_165 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c165
*+ bl_0_165 br_0_165 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c165
*+ bl_0_165 br_0_165 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c165
*+ bl_0_165 br_0_165 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c165
+ bl_0_165 br_0_165 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c166
+ bl_0_166 br_0_166 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c166
*+ bl_0_166 br_0_166 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c166
*+ bl_0_166 br_0_166 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c166
*+ bl_0_166 br_0_166 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c166
*+ bl_0_166 br_0_166 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c166
*+ bl_0_166 br_0_166 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c166
*+ bl_0_166 br_0_166 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c166
*+ bl_0_166 br_0_166 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c166
*+ bl_0_166 br_0_166 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c166
*+ bl_0_166 br_0_166 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c166
*+ bl_0_166 br_0_166 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c166
*+ bl_0_166 br_0_166 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c166
*+ bl_0_166 br_0_166 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c166
*+ bl_0_166 br_0_166 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c166
*+ bl_0_166 br_0_166 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c166
*+ bl_0_166 br_0_166 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c166
*+ bl_0_166 br_0_166 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c166
*+ bl_0_166 br_0_166 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c166
*+ bl_0_166 br_0_166 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c166
*+ bl_0_166 br_0_166 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c166
*+ bl_0_166 br_0_166 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c166
*+ bl_0_166 br_0_166 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c166
*+ bl_0_166 br_0_166 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c166
*+ bl_0_166 br_0_166 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c166
*+ bl_0_166 br_0_166 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c166
*+ bl_0_166 br_0_166 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c166
*+ bl_0_166 br_0_166 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c166
*+ bl_0_166 br_0_166 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c166
*+ bl_0_166 br_0_166 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c166
*+ bl_0_166 br_0_166 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c166
*+ bl_0_166 br_0_166 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c166
*+ bl_0_166 br_0_166 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c166
*+ bl_0_166 br_0_166 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c166
*+ bl_0_166 br_0_166 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c166
*+ bl_0_166 br_0_166 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c166
*+ bl_0_166 br_0_166 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c166
*+ bl_0_166 br_0_166 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c166
*+ bl_0_166 br_0_166 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c166
*+ bl_0_166 br_0_166 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c166
*+ bl_0_166 br_0_166 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c166
*+ bl_0_166 br_0_166 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c166
*+ bl_0_166 br_0_166 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c166
*+ bl_0_166 br_0_166 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c166
*+ bl_0_166 br_0_166 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c166
*+ bl_0_166 br_0_166 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c166
*+ bl_0_166 br_0_166 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c166
*+ bl_0_166 br_0_166 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c166
*+ bl_0_166 br_0_166 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c166
*+ bl_0_166 br_0_166 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c166
*+ bl_0_166 br_0_166 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c166
*+ bl_0_166 br_0_166 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c166
*+ bl_0_166 br_0_166 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c166
*+ bl_0_166 br_0_166 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c166
*+ bl_0_166 br_0_166 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c166
*+ bl_0_166 br_0_166 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c166
*+ bl_0_166 br_0_166 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c166
*+ bl_0_166 br_0_166 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c166
*+ bl_0_166 br_0_166 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c166
*+ bl_0_166 br_0_166 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c166
*+ bl_0_166 br_0_166 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c166
*+ bl_0_166 br_0_166 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c166
*+ bl_0_166 br_0_166 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c166
*+ bl_0_166 br_0_166 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c166
*+ bl_0_166 br_0_166 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c166
*+ bl_0_166 br_0_166 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c166
*+ bl_0_166 br_0_166 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c166
*+ bl_0_166 br_0_166 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c166
*+ bl_0_166 br_0_166 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c166
*+ bl_0_166 br_0_166 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c166
*+ bl_0_166 br_0_166 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c166
*+ bl_0_166 br_0_166 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c166
*+ bl_0_166 br_0_166 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c166
*+ bl_0_166 br_0_166 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c166
*+ bl_0_166 br_0_166 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c166
*+ bl_0_166 br_0_166 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c166
*+ bl_0_166 br_0_166 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c166
*+ bl_0_166 br_0_166 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c166
*+ bl_0_166 br_0_166 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c166
*+ bl_0_166 br_0_166 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c166
*+ bl_0_166 br_0_166 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c166
*+ bl_0_166 br_0_166 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c166
*+ bl_0_166 br_0_166 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c166
*+ bl_0_166 br_0_166 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c166
*+ bl_0_166 br_0_166 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c166
*+ bl_0_166 br_0_166 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c166
*+ bl_0_166 br_0_166 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c166
*+ bl_0_166 br_0_166 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c166
*+ bl_0_166 br_0_166 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c166
*+ bl_0_166 br_0_166 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c166
*+ bl_0_166 br_0_166 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c166
*+ bl_0_166 br_0_166 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c166
*+ bl_0_166 br_0_166 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c166
*+ bl_0_166 br_0_166 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c166
*+ bl_0_166 br_0_166 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c166
*+ bl_0_166 br_0_166 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c166
*+ bl_0_166 br_0_166 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c166
*+ bl_0_166 br_0_166 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c166
*+ bl_0_166 br_0_166 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c166
*+ bl_0_166 br_0_166 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c166
*+ bl_0_166 br_0_166 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c166
*+ bl_0_166 br_0_166 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c166
*+ bl_0_166 br_0_166 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c166
*+ bl_0_166 br_0_166 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c166
*+ bl_0_166 br_0_166 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c166
*+ bl_0_166 br_0_166 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c166
*+ bl_0_166 br_0_166 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c166
*+ bl_0_166 br_0_166 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c166
*+ bl_0_166 br_0_166 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c166
*+ bl_0_166 br_0_166 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c166
*+ bl_0_166 br_0_166 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c166
*+ bl_0_166 br_0_166 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c166
*+ bl_0_166 br_0_166 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c166
*+ bl_0_166 br_0_166 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c166
*+ bl_0_166 br_0_166 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c166
*+ bl_0_166 br_0_166 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c166
*+ bl_0_166 br_0_166 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c166
*+ bl_0_166 br_0_166 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c166
*+ bl_0_166 br_0_166 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c166
*+ bl_0_166 br_0_166 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c166
*+ bl_0_166 br_0_166 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c166
*+ bl_0_166 br_0_166 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c166
*+ bl_0_166 br_0_166 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c166
*+ bl_0_166 br_0_166 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c166
*+ bl_0_166 br_0_166 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c166
*+ bl_0_166 br_0_166 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c166
*+ bl_0_166 br_0_166 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c166
*+ bl_0_166 br_0_166 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c166
+ bl_0_166 br_0_166 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c167
+ bl_0_167 br_0_167 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c167
*+ bl_0_167 br_0_167 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c167
*+ bl_0_167 br_0_167 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c167
*+ bl_0_167 br_0_167 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c167
*+ bl_0_167 br_0_167 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c167
*+ bl_0_167 br_0_167 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c167
*+ bl_0_167 br_0_167 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c167
*+ bl_0_167 br_0_167 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c167
*+ bl_0_167 br_0_167 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c167
*+ bl_0_167 br_0_167 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c167
*+ bl_0_167 br_0_167 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c167
*+ bl_0_167 br_0_167 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c167
*+ bl_0_167 br_0_167 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c167
*+ bl_0_167 br_0_167 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c167
*+ bl_0_167 br_0_167 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c167
*+ bl_0_167 br_0_167 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c167
*+ bl_0_167 br_0_167 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c167
*+ bl_0_167 br_0_167 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c167
*+ bl_0_167 br_0_167 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c167
*+ bl_0_167 br_0_167 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c167
*+ bl_0_167 br_0_167 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c167
*+ bl_0_167 br_0_167 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c167
*+ bl_0_167 br_0_167 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c167
*+ bl_0_167 br_0_167 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c167
*+ bl_0_167 br_0_167 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c167
*+ bl_0_167 br_0_167 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c167
*+ bl_0_167 br_0_167 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c167
*+ bl_0_167 br_0_167 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c167
*+ bl_0_167 br_0_167 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c167
*+ bl_0_167 br_0_167 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c167
*+ bl_0_167 br_0_167 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c167
*+ bl_0_167 br_0_167 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c167
*+ bl_0_167 br_0_167 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c167
*+ bl_0_167 br_0_167 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c167
*+ bl_0_167 br_0_167 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c167
*+ bl_0_167 br_0_167 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c167
*+ bl_0_167 br_0_167 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c167
*+ bl_0_167 br_0_167 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c167
*+ bl_0_167 br_0_167 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c167
*+ bl_0_167 br_0_167 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c167
*+ bl_0_167 br_0_167 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c167
*+ bl_0_167 br_0_167 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c167
*+ bl_0_167 br_0_167 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c167
*+ bl_0_167 br_0_167 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c167
*+ bl_0_167 br_0_167 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c167
*+ bl_0_167 br_0_167 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c167
*+ bl_0_167 br_0_167 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c167
*+ bl_0_167 br_0_167 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c167
*+ bl_0_167 br_0_167 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c167
*+ bl_0_167 br_0_167 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c167
*+ bl_0_167 br_0_167 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c167
*+ bl_0_167 br_0_167 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c167
*+ bl_0_167 br_0_167 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c167
*+ bl_0_167 br_0_167 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c167
*+ bl_0_167 br_0_167 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c167
*+ bl_0_167 br_0_167 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c167
*+ bl_0_167 br_0_167 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c167
*+ bl_0_167 br_0_167 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c167
*+ bl_0_167 br_0_167 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c167
*+ bl_0_167 br_0_167 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c167
*+ bl_0_167 br_0_167 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c167
*+ bl_0_167 br_0_167 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c167
*+ bl_0_167 br_0_167 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c167
*+ bl_0_167 br_0_167 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c167
*+ bl_0_167 br_0_167 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c167
*+ bl_0_167 br_0_167 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c167
*+ bl_0_167 br_0_167 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c167
*+ bl_0_167 br_0_167 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c167
*+ bl_0_167 br_0_167 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c167
*+ bl_0_167 br_0_167 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c167
*+ bl_0_167 br_0_167 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c167
*+ bl_0_167 br_0_167 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c167
*+ bl_0_167 br_0_167 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c167
*+ bl_0_167 br_0_167 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c167
*+ bl_0_167 br_0_167 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c167
*+ bl_0_167 br_0_167 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c167
*+ bl_0_167 br_0_167 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c167
*+ bl_0_167 br_0_167 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c167
*+ bl_0_167 br_0_167 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c167
*+ bl_0_167 br_0_167 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c167
*+ bl_0_167 br_0_167 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c167
*+ bl_0_167 br_0_167 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c167
*+ bl_0_167 br_0_167 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c167
*+ bl_0_167 br_0_167 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c167
*+ bl_0_167 br_0_167 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c167
*+ bl_0_167 br_0_167 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c167
*+ bl_0_167 br_0_167 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c167
*+ bl_0_167 br_0_167 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c167
*+ bl_0_167 br_0_167 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c167
*+ bl_0_167 br_0_167 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c167
*+ bl_0_167 br_0_167 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c167
*+ bl_0_167 br_0_167 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c167
*+ bl_0_167 br_0_167 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c167
*+ bl_0_167 br_0_167 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c167
*+ bl_0_167 br_0_167 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c167
*+ bl_0_167 br_0_167 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c167
*+ bl_0_167 br_0_167 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c167
*+ bl_0_167 br_0_167 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c167
*+ bl_0_167 br_0_167 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c167
*+ bl_0_167 br_0_167 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c167
*+ bl_0_167 br_0_167 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c167
*+ bl_0_167 br_0_167 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c167
*+ bl_0_167 br_0_167 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c167
*+ bl_0_167 br_0_167 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c167
*+ bl_0_167 br_0_167 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c167
*+ bl_0_167 br_0_167 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c167
*+ bl_0_167 br_0_167 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c167
*+ bl_0_167 br_0_167 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c167
*+ bl_0_167 br_0_167 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c167
*+ bl_0_167 br_0_167 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c167
*+ bl_0_167 br_0_167 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c167
*+ bl_0_167 br_0_167 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c167
*+ bl_0_167 br_0_167 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c167
*+ bl_0_167 br_0_167 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c167
*+ bl_0_167 br_0_167 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c167
*+ bl_0_167 br_0_167 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c167
*+ bl_0_167 br_0_167 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c167
*+ bl_0_167 br_0_167 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c167
*+ bl_0_167 br_0_167 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c167
*+ bl_0_167 br_0_167 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c167
*+ bl_0_167 br_0_167 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c167
*+ bl_0_167 br_0_167 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c167
*+ bl_0_167 br_0_167 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c167
*+ bl_0_167 br_0_167 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c167
*+ bl_0_167 br_0_167 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c167
*+ bl_0_167 br_0_167 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c167
*+ bl_0_167 br_0_167 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c167
+ bl_0_167 br_0_167 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c168
+ bl_0_168 br_0_168 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c168
*+ bl_0_168 br_0_168 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c168
*+ bl_0_168 br_0_168 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c168
*+ bl_0_168 br_0_168 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c168
*+ bl_0_168 br_0_168 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c168
*+ bl_0_168 br_0_168 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c168
*+ bl_0_168 br_0_168 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c168
*+ bl_0_168 br_0_168 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c168
*+ bl_0_168 br_0_168 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c168
*+ bl_0_168 br_0_168 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c168
*+ bl_0_168 br_0_168 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c168
*+ bl_0_168 br_0_168 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c168
*+ bl_0_168 br_0_168 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c168
*+ bl_0_168 br_0_168 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c168
*+ bl_0_168 br_0_168 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c168
*+ bl_0_168 br_0_168 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c168
*+ bl_0_168 br_0_168 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c168
*+ bl_0_168 br_0_168 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c168
*+ bl_0_168 br_0_168 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c168
*+ bl_0_168 br_0_168 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c168
*+ bl_0_168 br_0_168 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c168
*+ bl_0_168 br_0_168 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c168
*+ bl_0_168 br_0_168 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c168
*+ bl_0_168 br_0_168 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c168
*+ bl_0_168 br_0_168 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c168
*+ bl_0_168 br_0_168 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c168
*+ bl_0_168 br_0_168 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c168
*+ bl_0_168 br_0_168 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c168
*+ bl_0_168 br_0_168 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c168
*+ bl_0_168 br_0_168 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c168
*+ bl_0_168 br_0_168 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c168
*+ bl_0_168 br_0_168 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c168
*+ bl_0_168 br_0_168 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c168
*+ bl_0_168 br_0_168 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c168
*+ bl_0_168 br_0_168 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c168
*+ bl_0_168 br_0_168 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c168
*+ bl_0_168 br_0_168 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c168
*+ bl_0_168 br_0_168 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c168
*+ bl_0_168 br_0_168 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c168
*+ bl_0_168 br_0_168 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c168
*+ bl_0_168 br_0_168 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c168
*+ bl_0_168 br_0_168 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c168
*+ bl_0_168 br_0_168 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c168
*+ bl_0_168 br_0_168 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c168
*+ bl_0_168 br_0_168 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c168
*+ bl_0_168 br_0_168 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c168
*+ bl_0_168 br_0_168 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c168
*+ bl_0_168 br_0_168 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c168
*+ bl_0_168 br_0_168 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c168
*+ bl_0_168 br_0_168 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c168
*+ bl_0_168 br_0_168 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c168
*+ bl_0_168 br_0_168 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c168
*+ bl_0_168 br_0_168 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c168
*+ bl_0_168 br_0_168 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c168
*+ bl_0_168 br_0_168 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c168
*+ bl_0_168 br_0_168 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c168
*+ bl_0_168 br_0_168 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c168
*+ bl_0_168 br_0_168 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c168
*+ bl_0_168 br_0_168 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c168
*+ bl_0_168 br_0_168 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c168
*+ bl_0_168 br_0_168 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c168
*+ bl_0_168 br_0_168 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c168
*+ bl_0_168 br_0_168 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c168
*+ bl_0_168 br_0_168 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c168
*+ bl_0_168 br_0_168 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c168
*+ bl_0_168 br_0_168 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c168
*+ bl_0_168 br_0_168 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c168
*+ bl_0_168 br_0_168 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c168
*+ bl_0_168 br_0_168 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c168
*+ bl_0_168 br_0_168 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c168
*+ bl_0_168 br_0_168 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c168
*+ bl_0_168 br_0_168 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c168
*+ bl_0_168 br_0_168 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c168
*+ bl_0_168 br_0_168 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c168
*+ bl_0_168 br_0_168 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c168
*+ bl_0_168 br_0_168 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c168
*+ bl_0_168 br_0_168 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c168
*+ bl_0_168 br_0_168 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c168
*+ bl_0_168 br_0_168 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c168
*+ bl_0_168 br_0_168 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c168
*+ bl_0_168 br_0_168 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c168
*+ bl_0_168 br_0_168 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c168
*+ bl_0_168 br_0_168 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c168
*+ bl_0_168 br_0_168 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c168
*+ bl_0_168 br_0_168 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c168
*+ bl_0_168 br_0_168 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c168
*+ bl_0_168 br_0_168 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c168
*+ bl_0_168 br_0_168 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c168
*+ bl_0_168 br_0_168 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c168
*+ bl_0_168 br_0_168 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c168
*+ bl_0_168 br_0_168 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c168
*+ bl_0_168 br_0_168 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c168
*+ bl_0_168 br_0_168 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c168
*+ bl_0_168 br_0_168 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c168
*+ bl_0_168 br_0_168 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c168
*+ bl_0_168 br_0_168 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c168
*+ bl_0_168 br_0_168 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c168
*+ bl_0_168 br_0_168 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c168
*+ bl_0_168 br_0_168 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c168
*+ bl_0_168 br_0_168 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c168
*+ bl_0_168 br_0_168 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c168
*+ bl_0_168 br_0_168 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c168
*+ bl_0_168 br_0_168 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c168
*+ bl_0_168 br_0_168 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c168
*+ bl_0_168 br_0_168 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c168
*+ bl_0_168 br_0_168 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c168
*+ bl_0_168 br_0_168 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c168
*+ bl_0_168 br_0_168 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c168
*+ bl_0_168 br_0_168 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c168
*+ bl_0_168 br_0_168 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c168
*+ bl_0_168 br_0_168 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c168
*+ bl_0_168 br_0_168 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c168
*+ bl_0_168 br_0_168 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c168
*+ bl_0_168 br_0_168 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c168
*+ bl_0_168 br_0_168 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c168
*+ bl_0_168 br_0_168 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c168
*+ bl_0_168 br_0_168 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c168
*+ bl_0_168 br_0_168 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c168
*+ bl_0_168 br_0_168 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c168
*+ bl_0_168 br_0_168 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c168
*+ bl_0_168 br_0_168 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c168
*+ bl_0_168 br_0_168 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c168
*+ bl_0_168 br_0_168 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c168
*+ bl_0_168 br_0_168 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c168
*+ bl_0_168 br_0_168 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c168
*+ bl_0_168 br_0_168 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c168
*+ bl_0_168 br_0_168 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c168
+ bl_0_168 br_0_168 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c169
+ bl_0_169 br_0_169 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c169
*+ bl_0_169 br_0_169 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c169
*+ bl_0_169 br_0_169 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c169
*+ bl_0_169 br_0_169 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c169
*+ bl_0_169 br_0_169 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c169
*+ bl_0_169 br_0_169 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c169
*+ bl_0_169 br_0_169 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c169
*+ bl_0_169 br_0_169 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c169
*+ bl_0_169 br_0_169 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c169
*+ bl_0_169 br_0_169 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c169
*+ bl_0_169 br_0_169 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c169
*+ bl_0_169 br_0_169 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c169
*+ bl_0_169 br_0_169 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c169
*+ bl_0_169 br_0_169 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c169
*+ bl_0_169 br_0_169 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c169
*+ bl_0_169 br_0_169 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c169
*+ bl_0_169 br_0_169 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c169
*+ bl_0_169 br_0_169 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c169
*+ bl_0_169 br_0_169 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c169
*+ bl_0_169 br_0_169 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c169
*+ bl_0_169 br_0_169 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c169
*+ bl_0_169 br_0_169 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c169
*+ bl_0_169 br_0_169 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c169
*+ bl_0_169 br_0_169 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c169
*+ bl_0_169 br_0_169 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c169
*+ bl_0_169 br_0_169 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c169
*+ bl_0_169 br_0_169 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c169
*+ bl_0_169 br_0_169 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c169
*+ bl_0_169 br_0_169 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c169
*+ bl_0_169 br_0_169 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c169
*+ bl_0_169 br_0_169 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c169
*+ bl_0_169 br_0_169 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c169
*+ bl_0_169 br_0_169 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c169
*+ bl_0_169 br_0_169 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c169
*+ bl_0_169 br_0_169 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c169
*+ bl_0_169 br_0_169 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c169
*+ bl_0_169 br_0_169 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c169
*+ bl_0_169 br_0_169 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c169
*+ bl_0_169 br_0_169 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c169
*+ bl_0_169 br_0_169 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c169
*+ bl_0_169 br_0_169 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c169
*+ bl_0_169 br_0_169 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c169
*+ bl_0_169 br_0_169 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c169
*+ bl_0_169 br_0_169 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c169
*+ bl_0_169 br_0_169 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c169
*+ bl_0_169 br_0_169 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c169
*+ bl_0_169 br_0_169 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c169
*+ bl_0_169 br_0_169 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c169
*+ bl_0_169 br_0_169 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c169
*+ bl_0_169 br_0_169 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c169
*+ bl_0_169 br_0_169 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c169
*+ bl_0_169 br_0_169 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c169
*+ bl_0_169 br_0_169 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c169
*+ bl_0_169 br_0_169 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c169
*+ bl_0_169 br_0_169 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c169
*+ bl_0_169 br_0_169 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c169
*+ bl_0_169 br_0_169 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c169
*+ bl_0_169 br_0_169 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c169
*+ bl_0_169 br_0_169 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c169
*+ bl_0_169 br_0_169 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c169
*+ bl_0_169 br_0_169 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c169
*+ bl_0_169 br_0_169 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c169
*+ bl_0_169 br_0_169 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c169
*+ bl_0_169 br_0_169 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c169
*+ bl_0_169 br_0_169 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c169
*+ bl_0_169 br_0_169 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c169
*+ bl_0_169 br_0_169 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c169
*+ bl_0_169 br_0_169 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c169
*+ bl_0_169 br_0_169 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c169
*+ bl_0_169 br_0_169 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c169
*+ bl_0_169 br_0_169 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c169
*+ bl_0_169 br_0_169 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c169
*+ bl_0_169 br_0_169 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c169
*+ bl_0_169 br_0_169 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c169
*+ bl_0_169 br_0_169 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c169
*+ bl_0_169 br_0_169 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c169
*+ bl_0_169 br_0_169 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c169
*+ bl_0_169 br_0_169 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c169
*+ bl_0_169 br_0_169 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c169
*+ bl_0_169 br_0_169 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c169
*+ bl_0_169 br_0_169 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c169
*+ bl_0_169 br_0_169 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c169
*+ bl_0_169 br_0_169 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c169
*+ bl_0_169 br_0_169 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c169
*+ bl_0_169 br_0_169 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c169
*+ bl_0_169 br_0_169 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c169
*+ bl_0_169 br_0_169 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c169
*+ bl_0_169 br_0_169 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c169
*+ bl_0_169 br_0_169 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c169
*+ bl_0_169 br_0_169 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c169
*+ bl_0_169 br_0_169 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c169
*+ bl_0_169 br_0_169 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c169
*+ bl_0_169 br_0_169 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c169
*+ bl_0_169 br_0_169 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c169
*+ bl_0_169 br_0_169 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c169
*+ bl_0_169 br_0_169 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c169
*+ bl_0_169 br_0_169 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c169
*+ bl_0_169 br_0_169 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c169
*+ bl_0_169 br_0_169 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c169
*+ bl_0_169 br_0_169 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c169
*+ bl_0_169 br_0_169 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c169
*+ bl_0_169 br_0_169 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c169
*+ bl_0_169 br_0_169 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c169
*+ bl_0_169 br_0_169 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c169
*+ bl_0_169 br_0_169 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c169
*+ bl_0_169 br_0_169 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c169
*+ bl_0_169 br_0_169 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c169
*+ bl_0_169 br_0_169 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c169
*+ bl_0_169 br_0_169 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c169
*+ bl_0_169 br_0_169 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c169
*+ bl_0_169 br_0_169 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c169
*+ bl_0_169 br_0_169 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c169
*+ bl_0_169 br_0_169 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c169
*+ bl_0_169 br_0_169 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c169
*+ bl_0_169 br_0_169 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c169
*+ bl_0_169 br_0_169 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c169
*+ bl_0_169 br_0_169 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c169
*+ bl_0_169 br_0_169 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c169
*+ bl_0_169 br_0_169 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c169
*+ bl_0_169 br_0_169 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c169
*+ bl_0_169 br_0_169 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c169
*+ bl_0_169 br_0_169 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c169
*+ bl_0_169 br_0_169 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c169
*+ bl_0_169 br_0_169 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c169
*+ bl_0_169 br_0_169 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c169
*+ bl_0_169 br_0_169 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c169
*+ bl_0_169 br_0_169 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c169
+ bl_0_169 br_0_169 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c170
+ bl_0_170 br_0_170 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c170
*+ bl_0_170 br_0_170 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c170
*+ bl_0_170 br_0_170 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c170
*+ bl_0_170 br_0_170 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c170
*+ bl_0_170 br_0_170 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c170
*+ bl_0_170 br_0_170 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c170
*+ bl_0_170 br_0_170 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c170
*+ bl_0_170 br_0_170 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c170
*+ bl_0_170 br_0_170 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c170
*+ bl_0_170 br_0_170 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c170
*+ bl_0_170 br_0_170 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c170
*+ bl_0_170 br_0_170 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c170
*+ bl_0_170 br_0_170 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c170
*+ bl_0_170 br_0_170 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c170
*+ bl_0_170 br_0_170 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c170
*+ bl_0_170 br_0_170 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c170
*+ bl_0_170 br_0_170 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c170
*+ bl_0_170 br_0_170 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c170
*+ bl_0_170 br_0_170 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c170
*+ bl_0_170 br_0_170 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c170
*+ bl_0_170 br_0_170 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c170
*+ bl_0_170 br_0_170 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c170
*+ bl_0_170 br_0_170 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c170
*+ bl_0_170 br_0_170 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c170
*+ bl_0_170 br_0_170 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c170
*+ bl_0_170 br_0_170 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c170
*+ bl_0_170 br_0_170 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c170
*+ bl_0_170 br_0_170 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c170
*+ bl_0_170 br_0_170 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c170
*+ bl_0_170 br_0_170 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c170
*+ bl_0_170 br_0_170 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c170
*+ bl_0_170 br_0_170 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c170
*+ bl_0_170 br_0_170 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c170
*+ bl_0_170 br_0_170 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c170
*+ bl_0_170 br_0_170 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c170
*+ bl_0_170 br_0_170 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c170
*+ bl_0_170 br_0_170 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c170
*+ bl_0_170 br_0_170 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c170
*+ bl_0_170 br_0_170 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c170
*+ bl_0_170 br_0_170 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c170
*+ bl_0_170 br_0_170 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c170
*+ bl_0_170 br_0_170 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c170
*+ bl_0_170 br_0_170 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c170
*+ bl_0_170 br_0_170 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c170
*+ bl_0_170 br_0_170 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c170
*+ bl_0_170 br_0_170 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c170
*+ bl_0_170 br_0_170 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c170
*+ bl_0_170 br_0_170 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c170
*+ bl_0_170 br_0_170 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c170
*+ bl_0_170 br_0_170 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c170
*+ bl_0_170 br_0_170 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c170
*+ bl_0_170 br_0_170 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c170
*+ bl_0_170 br_0_170 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c170
*+ bl_0_170 br_0_170 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c170
*+ bl_0_170 br_0_170 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c170
*+ bl_0_170 br_0_170 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c170
*+ bl_0_170 br_0_170 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c170
*+ bl_0_170 br_0_170 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c170
*+ bl_0_170 br_0_170 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c170
*+ bl_0_170 br_0_170 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c170
*+ bl_0_170 br_0_170 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c170
*+ bl_0_170 br_0_170 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c170
*+ bl_0_170 br_0_170 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c170
*+ bl_0_170 br_0_170 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c170
*+ bl_0_170 br_0_170 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c170
*+ bl_0_170 br_0_170 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c170
*+ bl_0_170 br_0_170 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c170
*+ bl_0_170 br_0_170 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c170
*+ bl_0_170 br_0_170 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c170
*+ bl_0_170 br_0_170 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c170
*+ bl_0_170 br_0_170 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c170
*+ bl_0_170 br_0_170 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c170
*+ bl_0_170 br_0_170 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c170
*+ bl_0_170 br_0_170 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c170
*+ bl_0_170 br_0_170 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c170
*+ bl_0_170 br_0_170 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c170
*+ bl_0_170 br_0_170 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c170
*+ bl_0_170 br_0_170 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c170
*+ bl_0_170 br_0_170 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c170
*+ bl_0_170 br_0_170 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c170
*+ bl_0_170 br_0_170 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c170
*+ bl_0_170 br_0_170 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c170
*+ bl_0_170 br_0_170 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c170
*+ bl_0_170 br_0_170 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c170
*+ bl_0_170 br_0_170 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c170
*+ bl_0_170 br_0_170 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c170
*+ bl_0_170 br_0_170 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c170
*+ bl_0_170 br_0_170 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c170
*+ bl_0_170 br_0_170 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c170
*+ bl_0_170 br_0_170 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c170
*+ bl_0_170 br_0_170 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c170
*+ bl_0_170 br_0_170 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c170
*+ bl_0_170 br_0_170 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c170
*+ bl_0_170 br_0_170 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c170
*+ bl_0_170 br_0_170 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c170
*+ bl_0_170 br_0_170 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c170
*+ bl_0_170 br_0_170 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c170
*+ bl_0_170 br_0_170 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c170
*+ bl_0_170 br_0_170 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c170
*+ bl_0_170 br_0_170 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c170
*+ bl_0_170 br_0_170 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c170
*+ bl_0_170 br_0_170 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c170
*+ bl_0_170 br_0_170 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c170
*+ bl_0_170 br_0_170 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c170
*+ bl_0_170 br_0_170 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c170
*+ bl_0_170 br_0_170 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c170
*+ bl_0_170 br_0_170 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c170
*+ bl_0_170 br_0_170 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c170
*+ bl_0_170 br_0_170 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c170
*+ bl_0_170 br_0_170 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c170
*+ bl_0_170 br_0_170 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c170
*+ bl_0_170 br_0_170 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c170
*+ bl_0_170 br_0_170 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c170
*+ bl_0_170 br_0_170 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c170
*+ bl_0_170 br_0_170 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c170
*+ bl_0_170 br_0_170 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c170
*+ bl_0_170 br_0_170 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c170
*+ bl_0_170 br_0_170 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c170
*+ bl_0_170 br_0_170 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c170
*+ bl_0_170 br_0_170 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c170
*+ bl_0_170 br_0_170 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c170
*+ bl_0_170 br_0_170 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c170
*+ bl_0_170 br_0_170 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c170
*+ bl_0_170 br_0_170 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c170
*+ bl_0_170 br_0_170 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c170
*+ bl_0_170 br_0_170 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c170
*+ bl_0_170 br_0_170 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c170
+ bl_0_170 br_0_170 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c171
+ bl_0_171 br_0_171 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c171
*+ bl_0_171 br_0_171 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c171
*+ bl_0_171 br_0_171 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c171
*+ bl_0_171 br_0_171 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c171
*+ bl_0_171 br_0_171 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c171
*+ bl_0_171 br_0_171 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c171
*+ bl_0_171 br_0_171 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c171
*+ bl_0_171 br_0_171 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c171
*+ bl_0_171 br_0_171 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c171
*+ bl_0_171 br_0_171 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c171
*+ bl_0_171 br_0_171 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c171
*+ bl_0_171 br_0_171 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c171
*+ bl_0_171 br_0_171 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c171
*+ bl_0_171 br_0_171 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c171
*+ bl_0_171 br_0_171 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c171
*+ bl_0_171 br_0_171 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c171
*+ bl_0_171 br_0_171 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c171
*+ bl_0_171 br_0_171 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c171
*+ bl_0_171 br_0_171 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c171
*+ bl_0_171 br_0_171 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c171
*+ bl_0_171 br_0_171 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c171
*+ bl_0_171 br_0_171 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c171
*+ bl_0_171 br_0_171 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c171
*+ bl_0_171 br_0_171 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c171
*+ bl_0_171 br_0_171 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c171
*+ bl_0_171 br_0_171 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c171
*+ bl_0_171 br_0_171 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c171
*+ bl_0_171 br_0_171 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c171
*+ bl_0_171 br_0_171 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c171
*+ bl_0_171 br_0_171 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c171
*+ bl_0_171 br_0_171 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c171
*+ bl_0_171 br_0_171 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c171
*+ bl_0_171 br_0_171 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c171
*+ bl_0_171 br_0_171 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c171
*+ bl_0_171 br_0_171 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c171
*+ bl_0_171 br_0_171 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c171
*+ bl_0_171 br_0_171 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c171
*+ bl_0_171 br_0_171 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c171
*+ bl_0_171 br_0_171 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c171
*+ bl_0_171 br_0_171 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c171
*+ bl_0_171 br_0_171 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c171
*+ bl_0_171 br_0_171 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c171
*+ bl_0_171 br_0_171 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c171
*+ bl_0_171 br_0_171 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c171
*+ bl_0_171 br_0_171 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c171
*+ bl_0_171 br_0_171 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c171
*+ bl_0_171 br_0_171 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c171
*+ bl_0_171 br_0_171 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c171
*+ bl_0_171 br_0_171 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c171
*+ bl_0_171 br_0_171 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c171
*+ bl_0_171 br_0_171 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c171
*+ bl_0_171 br_0_171 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c171
*+ bl_0_171 br_0_171 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c171
*+ bl_0_171 br_0_171 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c171
*+ bl_0_171 br_0_171 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c171
*+ bl_0_171 br_0_171 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c171
*+ bl_0_171 br_0_171 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c171
*+ bl_0_171 br_0_171 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c171
*+ bl_0_171 br_0_171 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c171
*+ bl_0_171 br_0_171 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c171
*+ bl_0_171 br_0_171 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c171
*+ bl_0_171 br_0_171 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c171
*+ bl_0_171 br_0_171 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c171
*+ bl_0_171 br_0_171 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c171
*+ bl_0_171 br_0_171 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c171
*+ bl_0_171 br_0_171 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c171
*+ bl_0_171 br_0_171 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c171
*+ bl_0_171 br_0_171 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c171
*+ bl_0_171 br_0_171 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c171
*+ bl_0_171 br_0_171 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c171
*+ bl_0_171 br_0_171 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c171
*+ bl_0_171 br_0_171 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c171
*+ bl_0_171 br_0_171 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c171
*+ bl_0_171 br_0_171 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c171
*+ bl_0_171 br_0_171 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c171
*+ bl_0_171 br_0_171 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c171
*+ bl_0_171 br_0_171 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c171
*+ bl_0_171 br_0_171 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c171
*+ bl_0_171 br_0_171 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c171
*+ bl_0_171 br_0_171 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c171
*+ bl_0_171 br_0_171 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c171
*+ bl_0_171 br_0_171 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c171
*+ bl_0_171 br_0_171 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c171
*+ bl_0_171 br_0_171 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c171
*+ bl_0_171 br_0_171 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c171
*+ bl_0_171 br_0_171 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c171
*+ bl_0_171 br_0_171 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c171
*+ bl_0_171 br_0_171 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c171
*+ bl_0_171 br_0_171 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c171
*+ bl_0_171 br_0_171 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c171
*+ bl_0_171 br_0_171 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c171
*+ bl_0_171 br_0_171 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c171
*+ bl_0_171 br_0_171 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c171
*+ bl_0_171 br_0_171 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c171
*+ bl_0_171 br_0_171 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c171
*+ bl_0_171 br_0_171 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c171
*+ bl_0_171 br_0_171 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c171
*+ bl_0_171 br_0_171 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c171
*+ bl_0_171 br_0_171 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c171
*+ bl_0_171 br_0_171 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c171
*+ bl_0_171 br_0_171 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c171
*+ bl_0_171 br_0_171 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c171
*+ bl_0_171 br_0_171 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c171
*+ bl_0_171 br_0_171 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c171
*+ bl_0_171 br_0_171 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c171
*+ bl_0_171 br_0_171 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c171
*+ bl_0_171 br_0_171 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c171
*+ bl_0_171 br_0_171 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c171
*+ bl_0_171 br_0_171 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c171
*+ bl_0_171 br_0_171 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c171
*+ bl_0_171 br_0_171 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c171
*+ bl_0_171 br_0_171 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c171
*+ bl_0_171 br_0_171 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c171
*+ bl_0_171 br_0_171 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c171
*+ bl_0_171 br_0_171 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c171
*+ bl_0_171 br_0_171 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c171
*+ bl_0_171 br_0_171 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c171
*+ bl_0_171 br_0_171 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c171
*+ bl_0_171 br_0_171 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c171
*+ bl_0_171 br_0_171 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c171
*+ bl_0_171 br_0_171 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c171
*+ bl_0_171 br_0_171 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c171
*+ bl_0_171 br_0_171 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c171
*+ bl_0_171 br_0_171 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c171
*+ bl_0_171 br_0_171 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c171
*+ bl_0_171 br_0_171 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c171
*+ bl_0_171 br_0_171 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c171
+ bl_0_171 br_0_171 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c172
+ bl_0_172 br_0_172 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c172
*+ bl_0_172 br_0_172 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c172
*+ bl_0_172 br_0_172 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c172
*+ bl_0_172 br_0_172 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c172
*+ bl_0_172 br_0_172 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c172
*+ bl_0_172 br_0_172 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c172
*+ bl_0_172 br_0_172 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c172
*+ bl_0_172 br_0_172 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c172
*+ bl_0_172 br_0_172 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c172
*+ bl_0_172 br_0_172 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c172
*+ bl_0_172 br_0_172 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c172
*+ bl_0_172 br_0_172 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c172
*+ bl_0_172 br_0_172 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c172
*+ bl_0_172 br_0_172 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c172
*+ bl_0_172 br_0_172 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c172
*+ bl_0_172 br_0_172 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c172
*+ bl_0_172 br_0_172 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c172
*+ bl_0_172 br_0_172 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c172
*+ bl_0_172 br_0_172 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c172
*+ bl_0_172 br_0_172 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c172
*+ bl_0_172 br_0_172 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c172
*+ bl_0_172 br_0_172 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c172
*+ bl_0_172 br_0_172 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c172
*+ bl_0_172 br_0_172 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c172
*+ bl_0_172 br_0_172 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c172
*+ bl_0_172 br_0_172 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c172
*+ bl_0_172 br_0_172 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c172
*+ bl_0_172 br_0_172 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c172
*+ bl_0_172 br_0_172 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c172
*+ bl_0_172 br_0_172 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c172
*+ bl_0_172 br_0_172 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c172
*+ bl_0_172 br_0_172 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c172
*+ bl_0_172 br_0_172 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c172
*+ bl_0_172 br_0_172 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c172
*+ bl_0_172 br_0_172 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c172
*+ bl_0_172 br_0_172 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c172
*+ bl_0_172 br_0_172 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c172
*+ bl_0_172 br_0_172 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c172
*+ bl_0_172 br_0_172 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c172
*+ bl_0_172 br_0_172 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c172
*+ bl_0_172 br_0_172 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c172
*+ bl_0_172 br_0_172 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c172
*+ bl_0_172 br_0_172 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c172
*+ bl_0_172 br_0_172 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c172
*+ bl_0_172 br_0_172 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c172
*+ bl_0_172 br_0_172 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c172
*+ bl_0_172 br_0_172 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c172
*+ bl_0_172 br_0_172 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c172
*+ bl_0_172 br_0_172 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c172
*+ bl_0_172 br_0_172 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c172
*+ bl_0_172 br_0_172 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c172
*+ bl_0_172 br_0_172 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c172
*+ bl_0_172 br_0_172 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c172
*+ bl_0_172 br_0_172 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c172
*+ bl_0_172 br_0_172 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c172
*+ bl_0_172 br_0_172 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c172
*+ bl_0_172 br_0_172 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c172
*+ bl_0_172 br_0_172 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c172
*+ bl_0_172 br_0_172 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c172
*+ bl_0_172 br_0_172 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c172
*+ bl_0_172 br_0_172 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c172
*+ bl_0_172 br_0_172 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c172
*+ bl_0_172 br_0_172 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c172
*+ bl_0_172 br_0_172 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c172
*+ bl_0_172 br_0_172 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c172
*+ bl_0_172 br_0_172 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c172
*+ bl_0_172 br_0_172 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c172
*+ bl_0_172 br_0_172 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c172
*+ bl_0_172 br_0_172 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c172
*+ bl_0_172 br_0_172 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c172
*+ bl_0_172 br_0_172 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c172
*+ bl_0_172 br_0_172 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c172
*+ bl_0_172 br_0_172 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c172
*+ bl_0_172 br_0_172 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c172
*+ bl_0_172 br_0_172 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c172
*+ bl_0_172 br_0_172 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c172
*+ bl_0_172 br_0_172 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c172
*+ bl_0_172 br_0_172 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c172
*+ bl_0_172 br_0_172 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c172
*+ bl_0_172 br_0_172 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c172
*+ bl_0_172 br_0_172 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c172
*+ bl_0_172 br_0_172 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c172
*+ bl_0_172 br_0_172 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c172
*+ bl_0_172 br_0_172 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c172
*+ bl_0_172 br_0_172 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c172
*+ bl_0_172 br_0_172 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c172
*+ bl_0_172 br_0_172 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c172
*+ bl_0_172 br_0_172 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c172
*+ bl_0_172 br_0_172 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c172
*+ bl_0_172 br_0_172 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c172
*+ bl_0_172 br_0_172 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c172
*+ bl_0_172 br_0_172 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c172
*+ bl_0_172 br_0_172 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c172
*+ bl_0_172 br_0_172 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c172
*+ bl_0_172 br_0_172 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c172
*+ bl_0_172 br_0_172 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c172
*+ bl_0_172 br_0_172 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c172
*+ bl_0_172 br_0_172 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c172
*+ bl_0_172 br_0_172 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c172
*+ bl_0_172 br_0_172 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c172
*+ bl_0_172 br_0_172 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c172
*+ bl_0_172 br_0_172 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c172
*+ bl_0_172 br_0_172 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c172
*+ bl_0_172 br_0_172 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c172
*+ bl_0_172 br_0_172 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c172
*+ bl_0_172 br_0_172 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c172
*+ bl_0_172 br_0_172 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c172
*+ bl_0_172 br_0_172 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c172
*+ bl_0_172 br_0_172 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c172
*+ bl_0_172 br_0_172 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c172
*+ bl_0_172 br_0_172 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c172
*+ bl_0_172 br_0_172 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c172
*+ bl_0_172 br_0_172 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c172
*+ bl_0_172 br_0_172 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c172
*+ bl_0_172 br_0_172 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c172
*+ bl_0_172 br_0_172 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c172
*+ bl_0_172 br_0_172 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c172
*+ bl_0_172 br_0_172 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c172
*+ bl_0_172 br_0_172 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c172
*+ bl_0_172 br_0_172 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c172
*+ bl_0_172 br_0_172 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c172
*+ bl_0_172 br_0_172 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c172
*+ bl_0_172 br_0_172 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c172
*+ bl_0_172 br_0_172 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c172
*+ bl_0_172 br_0_172 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c172
*+ bl_0_172 br_0_172 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c172
*+ bl_0_172 br_0_172 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c172
+ bl_0_172 br_0_172 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c173
+ bl_0_173 br_0_173 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c173
*+ bl_0_173 br_0_173 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c173
*+ bl_0_173 br_0_173 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c173
*+ bl_0_173 br_0_173 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c173
*+ bl_0_173 br_0_173 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c173
*+ bl_0_173 br_0_173 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c173
*+ bl_0_173 br_0_173 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c173
*+ bl_0_173 br_0_173 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c173
*+ bl_0_173 br_0_173 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c173
*+ bl_0_173 br_0_173 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c173
*+ bl_0_173 br_0_173 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c173
*+ bl_0_173 br_0_173 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c173
*+ bl_0_173 br_0_173 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c173
*+ bl_0_173 br_0_173 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c173
*+ bl_0_173 br_0_173 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c173
*+ bl_0_173 br_0_173 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c173
*+ bl_0_173 br_0_173 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c173
*+ bl_0_173 br_0_173 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c173
*+ bl_0_173 br_0_173 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c173
*+ bl_0_173 br_0_173 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c173
*+ bl_0_173 br_0_173 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c173
*+ bl_0_173 br_0_173 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c173
*+ bl_0_173 br_0_173 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c173
*+ bl_0_173 br_0_173 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c173
*+ bl_0_173 br_0_173 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c173
*+ bl_0_173 br_0_173 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c173
*+ bl_0_173 br_0_173 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c173
*+ bl_0_173 br_0_173 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c173
*+ bl_0_173 br_0_173 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c173
*+ bl_0_173 br_0_173 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c173
*+ bl_0_173 br_0_173 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c173
*+ bl_0_173 br_0_173 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c173
*+ bl_0_173 br_0_173 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c173
*+ bl_0_173 br_0_173 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c173
*+ bl_0_173 br_0_173 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c173
*+ bl_0_173 br_0_173 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c173
*+ bl_0_173 br_0_173 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c173
*+ bl_0_173 br_0_173 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c173
*+ bl_0_173 br_0_173 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c173
*+ bl_0_173 br_0_173 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c173
*+ bl_0_173 br_0_173 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c173
*+ bl_0_173 br_0_173 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c173
*+ bl_0_173 br_0_173 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c173
*+ bl_0_173 br_0_173 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c173
*+ bl_0_173 br_0_173 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c173
*+ bl_0_173 br_0_173 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c173
*+ bl_0_173 br_0_173 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c173
*+ bl_0_173 br_0_173 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c173
*+ bl_0_173 br_0_173 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c173
*+ bl_0_173 br_0_173 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c173
*+ bl_0_173 br_0_173 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c173
*+ bl_0_173 br_0_173 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c173
*+ bl_0_173 br_0_173 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c173
*+ bl_0_173 br_0_173 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c173
*+ bl_0_173 br_0_173 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c173
*+ bl_0_173 br_0_173 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c173
*+ bl_0_173 br_0_173 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c173
*+ bl_0_173 br_0_173 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c173
*+ bl_0_173 br_0_173 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c173
*+ bl_0_173 br_0_173 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c173
*+ bl_0_173 br_0_173 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c173
*+ bl_0_173 br_0_173 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c173
*+ bl_0_173 br_0_173 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c173
*+ bl_0_173 br_0_173 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c173
*+ bl_0_173 br_0_173 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c173
*+ bl_0_173 br_0_173 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c173
*+ bl_0_173 br_0_173 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c173
*+ bl_0_173 br_0_173 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c173
*+ bl_0_173 br_0_173 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c173
*+ bl_0_173 br_0_173 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c173
*+ bl_0_173 br_0_173 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c173
*+ bl_0_173 br_0_173 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c173
*+ bl_0_173 br_0_173 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c173
*+ bl_0_173 br_0_173 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c173
*+ bl_0_173 br_0_173 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c173
*+ bl_0_173 br_0_173 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c173
*+ bl_0_173 br_0_173 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c173
*+ bl_0_173 br_0_173 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c173
*+ bl_0_173 br_0_173 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c173
*+ bl_0_173 br_0_173 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c173
*+ bl_0_173 br_0_173 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c173
*+ bl_0_173 br_0_173 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c173
*+ bl_0_173 br_0_173 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c173
*+ bl_0_173 br_0_173 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c173
*+ bl_0_173 br_0_173 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c173
*+ bl_0_173 br_0_173 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c173
*+ bl_0_173 br_0_173 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c173
*+ bl_0_173 br_0_173 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c173
*+ bl_0_173 br_0_173 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c173
*+ bl_0_173 br_0_173 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c173
*+ bl_0_173 br_0_173 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c173
*+ bl_0_173 br_0_173 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c173
*+ bl_0_173 br_0_173 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c173
*+ bl_0_173 br_0_173 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c173
*+ bl_0_173 br_0_173 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c173
*+ bl_0_173 br_0_173 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c173
*+ bl_0_173 br_0_173 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c173
*+ bl_0_173 br_0_173 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c173
*+ bl_0_173 br_0_173 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c173
*+ bl_0_173 br_0_173 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c173
*+ bl_0_173 br_0_173 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c173
*+ bl_0_173 br_0_173 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c173
*+ bl_0_173 br_0_173 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c173
*+ bl_0_173 br_0_173 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c173
*+ bl_0_173 br_0_173 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c173
*+ bl_0_173 br_0_173 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c173
*+ bl_0_173 br_0_173 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c173
*+ bl_0_173 br_0_173 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c173
*+ bl_0_173 br_0_173 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c173
*+ bl_0_173 br_0_173 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c173
*+ bl_0_173 br_0_173 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c173
*+ bl_0_173 br_0_173 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c173
*+ bl_0_173 br_0_173 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c173
*+ bl_0_173 br_0_173 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c173
*+ bl_0_173 br_0_173 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c173
*+ bl_0_173 br_0_173 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c173
*+ bl_0_173 br_0_173 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c173
*+ bl_0_173 br_0_173 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c173
*+ bl_0_173 br_0_173 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c173
*+ bl_0_173 br_0_173 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c173
*+ bl_0_173 br_0_173 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c173
*+ bl_0_173 br_0_173 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c173
*+ bl_0_173 br_0_173 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c173
*+ bl_0_173 br_0_173 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c173
*+ bl_0_173 br_0_173 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c173
*+ bl_0_173 br_0_173 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c173
*+ bl_0_173 br_0_173 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c173
+ bl_0_173 br_0_173 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c174
+ bl_0_174 br_0_174 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c174
*+ bl_0_174 br_0_174 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c174
*+ bl_0_174 br_0_174 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c174
*+ bl_0_174 br_0_174 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c174
*+ bl_0_174 br_0_174 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c174
*+ bl_0_174 br_0_174 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c174
*+ bl_0_174 br_0_174 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c174
*+ bl_0_174 br_0_174 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c174
*+ bl_0_174 br_0_174 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c174
*+ bl_0_174 br_0_174 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c174
*+ bl_0_174 br_0_174 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c174
*+ bl_0_174 br_0_174 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c174
*+ bl_0_174 br_0_174 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c174
*+ bl_0_174 br_0_174 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c174
*+ bl_0_174 br_0_174 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c174
*+ bl_0_174 br_0_174 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c174
*+ bl_0_174 br_0_174 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c174
*+ bl_0_174 br_0_174 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c174
*+ bl_0_174 br_0_174 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c174
*+ bl_0_174 br_0_174 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c174
*+ bl_0_174 br_0_174 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c174
*+ bl_0_174 br_0_174 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c174
*+ bl_0_174 br_0_174 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c174
*+ bl_0_174 br_0_174 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c174
*+ bl_0_174 br_0_174 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c174
*+ bl_0_174 br_0_174 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c174
*+ bl_0_174 br_0_174 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c174
*+ bl_0_174 br_0_174 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c174
*+ bl_0_174 br_0_174 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c174
*+ bl_0_174 br_0_174 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c174
*+ bl_0_174 br_0_174 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c174
*+ bl_0_174 br_0_174 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c174
*+ bl_0_174 br_0_174 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c174
*+ bl_0_174 br_0_174 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c174
*+ bl_0_174 br_0_174 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c174
*+ bl_0_174 br_0_174 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c174
*+ bl_0_174 br_0_174 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c174
*+ bl_0_174 br_0_174 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c174
*+ bl_0_174 br_0_174 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c174
*+ bl_0_174 br_0_174 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c174
*+ bl_0_174 br_0_174 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c174
*+ bl_0_174 br_0_174 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c174
*+ bl_0_174 br_0_174 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c174
*+ bl_0_174 br_0_174 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c174
*+ bl_0_174 br_0_174 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c174
*+ bl_0_174 br_0_174 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c174
*+ bl_0_174 br_0_174 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c174
*+ bl_0_174 br_0_174 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c174
*+ bl_0_174 br_0_174 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c174
*+ bl_0_174 br_0_174 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c174
*+ bl_0_174 br_0_174 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c174
*+ bl_0_174 br_0_174 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c174
*+ bl_0_174 br_0_174 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c174
*+ bl_0_174 br_0_174 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c174
*+ bl_0_174 br_0_174 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c174
*+ bl_0_174 br_0_174 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c174
*+ bl_0_174 br_0_174 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c174
*+ bl_0_174 br_0_174 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c174
*+ bl_0_174 br_0_174 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c174
*+ bl_0_174 br_0_174 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c174
*+ bl_0_174 br_0_174 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c174
*+ bl_0_174 br_0_174 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c174
*+ bl_0_174 br_0_174 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c174
*+ bl_0_174 br_0_174 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c174
*+ bl_0_174 br_0_174 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c174
*+ bl_0_174 br_0_174 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c174
*+ bl_0_174 br_0_174 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c174
*+ bl_0_174 br_0_174 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c174
*+ bl_0_174 br_0_174 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c174
*+ bl_0_174 br_0_174 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c174
*+ bl_0_174 br_0_174 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c174
*+ bl_0_174 br_0_174 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c174
*+ bl_0_174 br_0_174 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c174
*+ bl_0_174 br_0_174 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c174
*+ bl_0_174 br_0_174 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c174
*+ bl_0_174 br_0_174 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c174
*+ bl_0_174 br_0_174 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c174
*+ bl_0_174 br_0_174 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c174
*+ bl_0_174 br_0_174 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c174
*+ bl_0_174 br_0_174 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c174
*+ bl_0_174 br_0_174 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c174
*+ bl_0_174 br_0_174 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c174
*+ bl_0_174 br_0_174 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c174
*+ bl_0_174 br_0_174 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c174
*+ bl_0_174 br_0_174 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c174
*+ bl_0_174 br_0_174 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c174
*+ bl_0_174 br_0_174 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c174
*+ bl_0_174 br_0_174 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c174
*+ bl_0_174 br_0_174 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c174
*+ bl_0_174 br_0_174 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c174
*+ bl_0_174 br_0_174 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c174
*+ bl_0_174 br_0_174 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c174
*+ bl_0_174 br_0_174 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c174
*+ bl_0_174 br_0_174 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c174
*+ bl_0_174 br_0_174 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c174
*+ bl_0_174 br_0_174 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c174
*+ bl_0_174 br_0_174 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c174
*+ bl_0_174 br_0_174 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c174
*+ bl_0_174 br_0_174 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c174
*+ bl_0_174 br_0_174 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c174
*+ bl_0_174 br_0_174 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c174
*+ bl_0_174 br_0_174 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c174
*+ bl_0_174 br_0_174 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c174
*+ bl_0_174 br_0_174 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c174
*+ bl_0_174 br_0_174 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c174
*+ bl_0_174 br_0_174 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c174
*+ bl_0_174 br_0_174 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c174
*+ bl_0_174 br_0_174 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c174
*+ bl_0_174 br_0_174 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c174
*+ bl_0_174 br_0_174 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c174
*+ bl_0_174 br_0_174 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c174
*+ bl_0_174 br_0_174 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c174
*+ bl_0_174 br_0_174 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c174
*+ bl_0_174 br_0_174 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c174
*+ bl_0_174 br_0_174 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c174
*+ bl_0_174 br_0_174 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c174
*+ bl_0_174 br_0_174 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c174
*+ bl_0_174 br_0_174 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c174
*+ bl_0_174 br_0_174 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c174
*+ bl_0_174 br_0_174 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c174
*+ bl_0_174 br_0_174 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c174
*+ bl_0_174 br_0_174 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c174
*+ bl_0_174 br_0_174 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c174
*+ bl_0_174 br_0_174 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c174
*+ bl_0_174 br_0_174 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c174
*+ bl_0_174 br_0_174 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c174
*+ bl_0_174 br_0_174 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c174
+ bl_0_174 br_0_174 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c175
+ bl_0_175 br_0_175 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c175
*+ bl_0_175 br_0_175 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c175
*+ bl_0_175 br_0_175 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c175
*+ bl_0_175 br_0_175 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c175
*+ bl_0_175 br_0_175 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c175
*+ bl_0_175 br_0_175 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c175
*+ bl_0_175 br_0_175 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c175
*+ bl_0_175 br_0_175 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c175
*+ bl_0_175 br_0_175 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c175
*+ bl_0_175 br_0_175 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c175
*+ bl_0_175 br_0_175 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c175
*+ bl_0_175 br_0_175 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c175
*+ bl_0_175 br_0_175 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c175
*+ bl_0_175 br_0_175 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c175
*+ bl_0_175 br_0_175 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c175
*+ bl_0_175 br_0_175 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c175
*+ bl_0_175 br_0_175 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c175
*+ bl_0_175 br_0_175 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c175
*+ bl_0_175 br_0_175 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c175
*+ bl_0_175 br_0_175 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c175
*+ bl_0_175 br_0_175 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c175
*+ bl_0_175 br_0_175 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c175
*+ bl_0_175 br_0_175 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c175
*+ bl_0_175 br_0_175 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c175
*+ bl_0_175 br_0_175 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c175
*+ bl_0_175 br_0_175 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c175
*+ bl_0_175 br_0_175 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c175
*+ bl_0_175 br_0_175 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c175
*+ bl_0_175 br_0_175 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c175
*+ bl_0_175 br_0_175 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c175
*+ bl_0_175 br_0_175 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c175
*+ bl_0_175 br_0_175 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c175
*+ bl_0_175 br_0_175 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c175
*+ bl_0_175 br_0_175 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c175
*+ bl_0_175 br_0_175 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c175
*+ bl_0_175 br_0_175 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c175
*+ bl_0_175 br_0_175 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c175
*+ bl_0_175 br_0_175 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c175
*+ bl_0_175 br_0_175 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c175
*+ bl_0_175 br_0_175 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c175
*+ bl_0_175 br_0_175 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c175
*+ bl_0_175 br_0_175 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c175
*+ bl_0_175 br_0_175 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c175
*+ bl_0_175 br_0_175 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c175
*+ bl_0_175 br_0_175 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c175
*+ bl_0_175 br_0_175 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c175
*+ bl_0_175 br_0_175 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c175
*+ bl_0_175 br_0_175 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c175
*+ bl_0_175 br_0_175 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c175
*+ bl_0_175 br_0_175 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c175
*+ bl_0_175 br_0_175 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c175
*+ bl_0_175 br_0_175 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c175
*+ bl_0_175 br_0_175 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c175
*+ bl_0_175 br_0_175 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c175
*+ bl_0_175 br_0_175 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c175
*+ bl_0_175 br_0_175 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c175
*+ bl_0_175 br_0_175 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c175
*+ bl_0_175 br_0_175 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c175
*+ bl_0_175 br_0_175 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c175
*+ bl_0_175 br_0_175 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c175
*+ bl_0_175 br_0_175 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c175
*+ bl_0_175 br_0_175 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c175
*+ bl_0_175 br_0_175 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c175
*+ bl_0_175 br_0_175 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c175
*+ bl_0_175 br_0_175 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c175
*+ bl_0_175 br_0_175 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c175
*+ bl_0_175 br_0_175 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c175
*+ bl_0_175 br_0_175 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c175
*+ bl_0_175 br_0_175 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c175
*+ bl_0_175 br_0_175 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c175
*+ bl_0_175 br_0_175 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c175
*+ bl_0_175 br_0_175 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c175
*+ bl_0_175 br_0_175 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c175
*+ bl_0_175 br_0_175 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c175
*+ bl_0_175 br_0_175 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c175
*+ bl_0_175 br_0_175 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c175
*+ bl_0_175 br_0_175 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c175
*+ bl_0_175 br_0_175 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c175
*+ bl_0_175 br_0_175 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c175
*+ bl_0_175 br_0_175 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c175
*+ bl_0_175 br_0_175 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c175
*+ bl_0_175 br_0_175 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c175
*+ bl_0_175 br_0_175 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c175
*+ bl_0_175 br_0_175 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c175
*+ bl_0_175 br_0_175 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c175
*+ bl_0_175 br_0_175 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c175
*+ bl_0_175 br_0_175 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c175
*+ bl_0_175 br_0_175 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c175
*+ bl_0_175 br_0_175 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c175
*+ bl_0_175 br_0_175 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c175
*+ bl_0_175 br_0_175 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c175
*+ bl_0_175 br_0_175 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c175
*+ bl_0_175 br_0_175 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c175
*+ bl_0_175 br_0_175 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c175
*+ bl_0_175 br_0_175 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c175
*+ bl_0_175 br_0_175 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c175
*+ bl_0_175 br_0_175 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c175
*+ bl_0_175 br_0_175 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c175
*+ bl_0_175 br_0_175 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c175
*+ bl_0_175 br_0_175 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c175
*+ bl_0_175 br_0_175 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c175
*+ bl_0_175 br_0_175 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c175
*+ bl_0_175 br_0_175 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c175
*+ bl_0_175 br_0_175 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c175
*+ bl_0_175 br_0_175 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c175
*+ bl_0_175 br_0_175 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c175
*+ bl_0_175 br_0_175 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c175
*+ bl_0_175 br_0_175 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c175
*+ bl_0_175 br_0_175 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c175
*+ bl_0_175 br_0_175 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c175
*+ bl_0_175 br_0_175 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c175
*+ bl_0_175 br_0_175 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c175
*+ bl_0_175 br_0_175 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c175
*+ bl_0_175 br_0_175 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c175
*+ bl_0_175 br_0_175 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c175
*+ bl_0_175 br_0_175 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c175
*+ bl_0_175 br_0_175 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c175
*+ bl_0_175 br_0_175 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c175
*+ bl_0_175 br_0_175 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c175
*+ bl_0_175 br_0_175 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c175
*+ bl_0_175 br_0_175 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c175
*+ bl_0_175 br_0_175 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c175
*+ bl_0_175 br_0_175 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c175
*+ bl_0_175 br_0_175 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c175
*+ bl_0_175 br_0_175 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c175
*+ bl_0_175 br_0_175 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c175
*+ bl_0_175 br_0_175 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c175
+ bl_0_175 br_0_175 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c176
+ bl_0_176 br_0_176 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c176
*+ bl_0_176 br_0_176 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c176
*+ bl_0_176 br_0_176 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c176
*+ bl_0_176 br_0_176 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c176
*+ bl_0_176 br_0_176 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c176
*+ bl_0_176 br_0_176 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c176
*+ bl_0_176 br_0_176 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c176
*+ bl_0_176 br_0_176 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c176
*+ bl_0_176 br_0_176 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c176
*+ bl_0_176 br_0_176 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c176
*+ bl_0_176 br_0_176 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c176
*+ bl_0_176 br_0_176 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c176
*+ bl_0_176 br_0_176 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c176
*+ bl_0_176 br_0_176 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c176
*+ bl_0_176 br_0_176 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c176
*+ bl_0_176 br_0_176 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c176
*+ bl_0_176 br_0_176 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c176
*+ bl_0_176 br_0_176 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c176
*+ bl_0_176 br_0_176 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c176
*+ bl_0_176 br_0_176 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c176
*+ bl_0_176 br_0_176 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c176
*+ bl_0_176 br_0_176 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c176
*+ bl_0_176 br_0_176 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c176
*+ bl_0_176 br_0_176 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c176
*+ bl_0_176 br_0_176 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c176
*+ bl_0_176 br_0_176 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c176
*+ bl_0_176 br_0_176 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c176
*+ bl_0_176 br_0_176 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c176
*+ bl_0_176 br_0_176 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c176
*+ bl_0_176 br_0_176 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c176
*+ bl_0_176 br_0_176 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c176
*+ bl_0_176 br_0_176 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c176
*+ bl_0_176 br_0_176 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c176
*+ bl_0_176 br_0_176 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c176
*+ bl_0_176 br_0_176 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c176
*+ bl_0_176 br_0_176 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c176
*+ bl_0_176 br_0_176 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c176
*+ bl_0_176 br_0_176 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c176
*+ bl_0_176 br_0_176 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c176
*+ bl_0_176 br_0_176 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c176
*+ bl_0_176 br_0_176 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c176
*+ bl_0_176 br_0_176 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c176
*+ bl_0_176 br_0_176 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c176
*+ bl_0_176 br_0_176 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c176
*+ bl_0_176 br_0_176 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c176
*+ bl_0_176 br_0_176 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c176
*+ bl_0_176 br_0_176 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c176
*+ bl_0_176 br_0_176 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c176
*+ bl_0_176 br_0_176 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c176
*+ bl_0_176 br_0_176 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c176
*+ bl_0_176 br_0_176 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c176
*+ bl_0_176 br_0_176 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c176
*+ bl_0_176 br_0_176 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c176
*+ bl_0_176 br_0_176 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c176
*+ bl_0_176 br_0_176 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c176
*+ bl_0_176 br_0_176 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c176
*+ bl_0_176 br_0_176 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c176
*+ bl_0_176 br_0_176 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c176
*+ bl_0_176 br_0_176 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c176
*+ bl_0_176 br_0_176 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c176
*+ bl_0_176 br_0_176 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c176
*+ bl_0_176 br_0_176 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c176
*+ bl_0_176 br_0_176 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c176
*+ bl_0_176 br_0_176 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c176
*+ bl_0_176 br_0_176 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c176
*+ bl_0_176 br_0_176 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c176
*+ bl_0_176 br_0_176 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c176
*+ bl_0_176 br_0_176 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c176
*+ bl_0_176 br_0_176 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c176
*+ bl_0_176 br_0_176 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c176
*+ bl_0_176 br_0_176 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c176
*+ bl_0_176 br_0_176 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c176
*+ bl_0_176 br_0_176 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c176
*+ bl_0_176 br_0_176 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c176
*+ bl_0_176 br_0_176 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c176
*+ bl_0_176 br_0_176 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c176
*+ bl_0_176 br_0_176 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c176
*+ bl_0_176 br_0_176 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c176
*+ bl_0_176 br_0_176 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c176
*+ bl_0_176 br_0_176 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c176
*+ bl_0_176 br_0_176 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c176
*+ bl_0_176 br_0_176 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c176
*+ bl_0_176 br_0_176 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c176
*+ bl_0_176 br_0_176 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c176
*+ bl_0_176 br_0_176 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c176
*+ bl_0_176 br_0_176 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c176
*+ bl_0_176 br_0_176 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c176
*+ bl_0_176 br_0_176 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c176
*+ bl_0_176 br_0_176 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c176
*+ bl_0_176 br_0_176 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c176
*+ bl_0_176 br_0_176 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c176
*+ bl_0_176 br_0_176 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c176
*+ bl_0_176 br_0_176 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c176
*+ bl_0_176 br_0_176 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c176
*+ bl_0_176 br_0_176 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c176
*+ bl_0_176 br_0_176 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c176
*+ bl_0_176 br_0_176 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c176
*+ bl_0_176 br_0_176 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c176
*+ bl_0_176 br_0_176 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c176
*+ bl_0_176 br_0_176 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c176
*+ bl_0_176 br_0_176 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c176
*+ bl_0_176 br_0_176 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c176
*+ bl_0_176 br_0_176 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c176
*+ bl_0_176 br_0_176 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c176
*+ bl_0_176 br_0_176 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c176
*+ bl_0_176 br_0_176 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c176
*+ bl_0_176 br_0_176 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c176
*+ bl_0_176 br_0_176 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c176
*+ bl_0_176 br_0_176 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c176
*+ bl_0_176 br_0_176 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c176
*+ bl_0_176 br_0_176 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c176
*+ bl_0_176 br_0_176 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c176
*+ bl_0_176 br_0_176 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c176
*+ bl_0_176 br_0_176 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c176
*+ bl_0_176 br_0_176 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c176
*+ bl_0_176 br_0_176 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c176
*+ bl_0_176 br_0_176 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c176
*+ bl_0_176 br_0_176 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c176
*+ bl_0_176 br_0_176 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c176
*+ bl_0_176 br_0_176 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c176
*+ bl_0_176 br_0_176 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c176
*+ bl_0_176 br_0_176 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c176
*+ bl_0_176 br_0_176 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c176
*+ bl_0_176 br_0_176 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c176
*+ bl_0_176 br_0_176 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c176
*+ bl_0_176 br_0_176 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c176
*+ bl_0_176 br_0_176 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c176
+ bl_0_176 br_0_176 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c177
+ bl_0_177 br_0_177 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c177
*+ bl_0_177 br_0_177 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c177
*+ bl_0_177 br_0_177 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c177
*+ bl_0_177 br_0_177 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c177
*+ bl_0_177 br_0_177 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c177
*+ bl_0_177 br_0_177 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c177
*+ bl_0_177 br_0_177 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c177
*+ bl_0_177 br_0_177 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c177
*+ bl_0_177 br_0_177 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c177
*+ bl_0_177 br_0_177 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c177
*+ bl_0_177 br_0_177 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c177
*+ bl_0_177 br_0_177 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c177
*+ bl_0_177 br_0_177 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c177
*+ bl_0_177 br_0_177 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c177
*+ bl_0_177 br_0_177 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c177
*+ bl_0_177 br_0_177 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c177
*+ bl_0_177 br_0_177 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c177
*+ bl_0_177 br_0_177 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c177
*+ bl_0_177 br_0_177 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c177
*+ bl_0_177 br_0_177 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c177
*+ bl_0_177 br_0_177 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c177
*+ bl_0_177 br_0_177 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c177
*+ bl_0_177 br_0_177 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c177
*+ bl_0_177 br_0_177 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c177
*+ bl_0_177 br_0_177 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c177
*+ bl_0_177 br_0_177 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c177
*+ bl_0_177 br_0_177 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c177
*+ bl_0_177 br_0_177 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c177
*+ bl_0_177 br_0_177 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c177
*+ bl_0_177 br_0_177 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c177
*+ bl_0_177 br_0_177 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c177
*+ bl_0_177 br_0_177 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c177
*+ bl_0_177 br_0_177 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c177
*+ bl_0_177 br_0_177 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c177
*+ bl_0_177 br_0_177 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c177
*+ bl_0_177 br_0_177 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c177
*+ bl_0_177 br_0_177 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c177
*+ bl_0_177 br_0_177 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c177
*+ bl_0_177 br_0_177 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c177
*+ bl_0_177 br_0_177 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c177
*+ bl_0_177 br_0_177 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c177
*+ bl_0_177 br_0_177 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c177
*+ bl_0_177 br_0_177 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c177
*+ bl_0_177 br_0_177 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c177
*+ bl_0_177 br_0_177 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c177
*+ bl_0_177 br_0_177 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c177
*+ bl_0_177 br_0_177 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c177
*+ bl_0_177 br_0_177 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c177
*+ bl_0_177 br_0_177 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c177
*+ bl_0_177 br_0_177 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c177
*+ bl_0_177 br_0_177 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c177
*+ bl_0_177 br_0_177 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c177
*+ bl_0_177 br_0_177 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c177
*+ bl_0_177 br_0_177 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c177
*+ bl_0_177 br_0_177 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c177
*+ bl_0_177 br_0_177 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c177
*+ bl_0_177 br_0_177 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c177
*+ bl_0_177 br_0_177 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c177
*+ bl_0_177 br_0_177 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c177
*+ bl_0_177 br_0_177 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c177
*+ bl_0_177 br_0_177 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c177
*+ bl_0_177 br_0_177 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c177
*+ bl_0_177 br_0_177 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c177
*+ bl_0_177 br_0_177 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c177
*+ bl_0_177 br_0_177 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c177
*+ bl_0_177 br_0_177 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c177
*+ bl_0_177 br_0_177 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c177
*+ bl_0_177 br_0_177 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c177
*+ bl_0_177 br_0_177 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c177
*+ bl_0_177 br_0_177 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c177
*+ bl_0_177 br_0_177 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c177
*+ bl_0_177 br_0_177 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c177
*+ bl_0_177 br_0_177 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c177
*+ bl_0_177 br_0_177 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c177
*+ bl_0_177 br_0_177 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c177
*+ bl_0_177 br_0_177 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c177
*+ bl_0_177 br_0_177 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c177
*+ bl_0_177 br_0_177 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c177
*+ bl_0_177 br_0_177 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c177
*+ bl_0_177 br_0_177 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c177
*+ bl_0_177 br_0_177 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c177
*+ bl_0_177 br_0_177 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c177
*+ bl_0_177 br_0_177 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c177
*+ bl_0_177 br_0_177 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c177
*+ bl_0_177 br_0_177 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c177
*+ bl_0_177 br_0_177 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c177
*+ bl_0_177 br_0_177 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c177
*+ bl_0_177 br_0_177 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c177
*+ bl_0_177 br_0_177 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c177
*+ bl_0_177 br_0_177 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c177
*+ bl_0_177 br_0_177 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c177
*+ bl_0_177 br_0_177 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c177
*+ bl_0_177 br_0_177 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c177
*+ bl_0_177 br_0_177 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c177
*+ bl_0_177 br_0_177 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c177
*+ bl_0_177 br_0_177 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c177
*+ bl_0_177 br_0_177 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c177
*+ bl_0_177 br_0_177 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c177
*+ bl_0_177 br_0_177 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c177
*+ bl_0_177 br_0_177 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c177
*+ bl_0_177 br_0_177 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c177
*+ bl_0_177 br_0_177 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c177
*+ bl_0_177 br_0_177 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c177
*+ bl_0_177 br_0_177 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c177
*+ bl_0_177 br_0_177 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c177
*+ bl_0_177 br_0_177 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c177
*+ bl_0_177 br_0_177 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c177
*+ bl_0_177 br_0_177 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c177
*+ bl_0_177 br_0_177 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c177
*+ bl_0_177 br_0_177 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c177
*+ bl_0_177 br_0_177 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c177
*+ bl_0_177 br_0_177 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c177
*+ bl_0_177 br_0_177 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c177
*+ bl_0_177 br_0_177 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c177
*+ bl_0_177 br_0_177 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c177
*+ bl_0_177 br_0_177 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c177
*+ bl_0_177 br_0_177 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c177
*+ bl_0_177 br_0_177 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c177
*+ bl_0_177 br_0_177 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c177
*+ bl_0_177 br_0_177 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c177
*+ bl_0_177 br_0_177 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c177
*+ bl_0_177 br_0_177 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c177
*+ bl_0_177 br_0_177 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c177
*+ bl_0_177 br_0_177 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c177
*+ bl_0_177 br_0_177 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c177
*+ bl_0_177 br_0_177 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c177
*+ bl_0_177 br_0_177 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c177
+ bl_0_177 br_0_177 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c178
+ bl_0_178 br_0_178 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c178
*+ bl_0_178 br_0_178 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c178
*+ bl_0_178 br_0_178 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c178
*+ bl_0_178 br_0_178 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c178
*+ bl_0_178 br_0_178 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c178
*+ bl_0_178 br_0_178 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c178
*+ bl_0_178 br_0_178 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c178
*+ bl_0_178 br_0_178 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c178
*+ bl_0_178 br_0_178 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c178
*+ bl_0_178 br_0_178 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c178
*+ bl_0_178 br_0_178 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c178
*+ bl_0_178 br_0_178 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c178
*+ bl_0_178 br_0_178 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c178
*+ bl_0_178 br_0_178 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c178
*+ bl_0_178 br_0_178 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c178
*+ bl_0_178 br_0_178 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c178
*+ bl_0_178 br_0_178 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c178
*+ bl_0_178 br_0_178 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c178
*+ bl_0_178 br_0_178 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c178
*+ bl_0_178 br_0_178 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c178
*+ bl_0_178 br_0_178 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c178
*+ bl_0_178 br_0_178 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c178
*+ bl_0_178 br_0_178 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c178
*+ bl_0_178 br_0_178 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c178
*+ bl_0_178 br_0_178 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c178
*+ bl_0_178 br_0_178 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c178
*+ bl_0_178 br_0_178 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c178
*+ bl_0_178 br_0_178 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c178
*+ bl_0_178 br_0_178 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c178
*+ bl_0_178 br_0_178 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c178
*+ bl_0_178 br_0_178 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c178
*+ bl_0_178 br_0_178 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c178
*+ bl_0_178 br_0_178 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c178
*+ bl_0_178 br_0_178 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c178
*+ bl_0_178 br_0_178 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c178
*+ bl_0_178 br_0_178 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c178
*+ bl_0_178 br_0_178 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c178
*+ bl_0_178 br_0_178 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c178
*+ bl_0_178 br_0_178 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c178
*+ bl_0_178 br_0_178 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c178
*+ bl_0_178 br_0_178 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c178
*+ bl_0_178 br_0_178 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c178
*+ bl_0_178 br_0_178 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c178
*+ bl_0_178 br_0_178 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c178
*+ bl_0_178 br_0_178 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c178
*+ bl_0_178 br_0_178 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c178
*+ bl_0_178 br_0_178 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c178
*+ bl_0_178 br_0_178 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c178
*+ bl_0_178 br_0_178 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c178
*+ bl_0_178 br_0_178 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c178
*+ bl_0_178 br_0_178 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c178
*+ bl_0_178 br_0_178 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c178
*+ bl_0_178 br_0_178 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c178
*+ bl_0_178 br_0_178 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c178
*+ bl_0_178 br_0_178 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c178
*+ bl_0_178 br_0_178 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c178
*+ bl_0_178 br_0_178 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c178
*+ bl_0_178 br_0_178 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c178
*+ bl_0_178 br_0_178 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c178
*+ bl_0_178 br_0_178 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c178
*+ bl_0_178 br_0_178 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c178
*+ bl_0_178 br_0_178 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c178
*+ bl_0_178 br_0_178 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c178
*+ bl_0_178 br_0_178 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c178
*+ bl_0_178 br_0_178 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c178
*+ bl_0_178 br_0_178 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c178
*+ bl_0_178 br_0_178 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c178
*+ bl_0_178 br_0_178 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c178
*+ bl_0_178 br_0_178 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c178
*+ bl_0_178 br_0_178 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c178
*+ bl_0_178 br_0_178 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c178
*+ bl_0_178 br_0_178 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c178
*+ bl_0_178 br_0_178 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c178
*+ bl_0_178 br_0_178 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c178
*+ bl_0_178 br_0_178 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c178
*+ bl_0_178 br_0_178 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c178
*+ bl_0_178 br_0_178 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c178
*+ bl_0_178 br_0_178 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c178
*+ bl_0_178 br_0_178 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c178
*+ bl_0_178 br_0_178 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c178
*+ bl_0_178 br_0_178 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c178
*+ bl_0_178 br_0_178 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c178
*+ bl_0_178 br_0_178 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c178
*+ bl_0_178 br_0_178 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c178
*+ bl_0_178 br_0_178 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c178
*+ bl_0_178 br_0_178 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c178
*+ bl_0_178 br_0_178 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c178
*+ bl_0_178 br_0_178 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c178
*+ bl_0_178 br_0_178 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c178
*+ bl_0_178 br_0_178 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c178
*+ bl_0_178 br_0_178 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c178
*+ bl_0_178 br_0_178 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c178
*+ bl_0_178 br_0_178 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c178
*+ bl_0_178 br_0_178 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c178
*+ bl_0_178 br_0_178 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c178
*+ bl_0_178 br_0_178 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c178
*+ bl_0_178 br_0_178 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c178
*+ bl_0_178 br_0_178 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c178
*+ bl_0_178 br_0_178 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c178
*+ bl_0_178 br_0_178 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c178
*+ bl_0_178 br_0_178 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c178
*+ bl_0_178 br_0_178 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c178
*+ bl_0_178 br_0_178 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c178
*+ bl_0_178 br_0_178 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c178
*+ bl_0_178 br_0_178 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c178
*+ bl_0_178 br_0_178 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c178
*+ bl_0_178 br_0_178 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c178
*+ bl_0_178 br_0_178 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c178
*+ bl_0_178 br_0_178 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c178
*+ bl_0_178 br_0_178 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c178
*+ bl_0_178 br_0_178 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c178
*+ bl_0_178 br_0_178 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c178
*+ bl_0_178 br_0_178 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c178
*+ bl_0_178 br_0_178 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c178
*+ bl_0_178 br_0_178 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c178
*+ bl_0_178 br_0_178 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c178
*+ bl_0_178 br_0_178 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c178
*+ bl_0_178 br_0_178 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c178
*+ bl_0_178 br_0_178 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c178
*+ bl_0_178 br_0_178 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c178
*+ bl_0_178 br_0_178 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c178
*+ bl_0_178 br_0_178 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c178
*+ bl_0_178 br_0_178 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c178
*+ bl_0_178 br_0_178 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c178
*+ bl_0_178 br_0_178 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c178
*+ bl_0_178 br_0_178 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c178
*+ bl_0_178 br_0_178 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c178
+ bl_0_178 br_0_178 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c179
+ bl_0_179 br_0_179 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c179
*+ bl_0_179 br_0_179 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c179
*+ bl_0_179 br_0_179 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c179
*+ bl_0_179 br_0_179 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c179
*+ bl_0_179 br_0_179 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c179
*+ bl_0_179 br_0_179 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c179
*+ bl_0_179 br_0_179 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c179
*+ bl_0_179 br_0_179 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c179
*+ bl_0_179 br_0_179 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c179
*+ bl_0_179 br_0_179 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c179
*+ bl_0_179 br_0_179 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c179
*+ bl_0_179 br_0_179 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c179
*+ bl_0_179 br_0_179 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c179
*+ bl_0_179 br_0_179 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c179
*+ bl_0_179 br_0_179 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c179
*+ bl_0_179 br_0_179 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c179
*+ bl_0_179 br_0_179 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c179
*+ bl_0_179 br_0_179 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c179
*+ bl_0_179 br_0_179 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c179
*+ bl_0_179 br_0_179 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c179
*+ bl_0_179 br_0_179 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c179
*+ bl_0_179 br_0_179 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c179
*+ bl_0_179 br_0_179 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c179
*+ bl_0_179 br_0_179 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c179
*+ bl_0_179 br_0_179 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c179
*+ bl_0_179 br_0_179 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c179
*+ bl_0_179 br_0_179 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c179
*+ bl_0_179 br_0_179 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c179
*+ bl_0_179 br_0_179 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c179
*+ bl_0_179 br_0_179 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c179
*+ bl_0_179 br_0_179 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c179
*+ bl_0_179 br_0_179 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c179
*+ bl_0_179 br_0_179 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c179
*+ bl_0_179 br_0_179 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c179
*+ bl_0_179 br_0_179 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c179
*+ bl_0_179 br_0_179 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c179
*+ bl_0_179 br_0_179 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c179
*+ bl_0_179 br_0_179 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c179
*+ bl_0_179 br_0_179 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c179
*+ bl_0_179 br_0_179 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c179
*+ bl_0_179 br_0_179 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c179
*+ bl_0_179 br_0_179 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c179
*+ bl_0_179 br_0_179 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c179
*+ bl_0_179 br_0_179 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c179
*+ bl_0_179 br_0_179 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c179
*+ bl_0_179 br_0_179 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c179
*+ bl_0_179 br_0_179 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c179
*+ bl_0_179 br_0_179 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c179
*+ bl_0_179 br_0_179 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c179
*+ bl_0_179 br_0_179 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c179
*+ bl_0_179 br_0_179 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c179
*+ bl_0_179 br_0_179 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c179
*+ bl_0_179 br_0_179 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c179
*+ bl_0_179 br_0_179 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c179
*+ bl_0_179 br_0_179 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c179
*+ bl_0_179 br_0_179 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c179
*+ bl_0_179 br_0_179 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c179
*+ bl_0_179 br_0_179 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c179
*+ bl_0_179 br_0_179 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c179
*+ bl_0_179 br_0_179 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c179
*+ bl_0_179 br_0_179 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c179
*+ bl_0_179 br_0_179 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c179
*+ bl_0_179 br_0_179 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c179
*+ bl_0_179 br_0_179 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c179
*+ bl_0_179 br_0_179 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c179
*+ bl_0_179 br_0_179 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c179
*+ bl_0_179 br_0_179 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c179
*+ bl_0_179 br_0_179 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c179
*+ bl_0_179 br_0_179 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c179
*+ bl_0_179 br_0_179 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c179
*+ bl_0_179 br_0_179 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c179
*+ bl_0_179 br_0_179 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c179
*+ bl_0_179 br_0_179 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c179
*+ bl_0_179 br_0_179 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c179
*+ bl_0_179 br_0_179 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c179
*+ bl_0_179 br_0_179 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c179
*+ bl_0_179 br_0_179 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c179
*+ bl_0_179 br_0_179 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c179
*+ bl_0_179 br_0_179 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c179
*+ bl_0_179 br_0_179 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c179
*+ bl_0_179 br_0_179 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c179
*+ bl_0_179 br_0_179 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c179
*+ bl_0_179 br_0_179 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c179
*+ bl_0_179 br_0_179 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c179
*+ bl_0_179 br_0_179 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c179
*+ bl_0_179 br_0_179 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c179
*+ bl_0_179 br_0_179 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c179
*+ bl_0_179 br_0_179 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c179
*+ bl_0_179 br_0_179 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c179
*+ bl_0_179 br_0_179 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c179
*+ bl_0_179 br_0_179 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c179
*+ bl_0_179 br_0_179 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c179
*+ bl_0_179 br_0_179 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c179
*+ bl_0_179 br_0_179 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c179
*+ bl_0_179 br_0_179 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c179
*+ bl_0_179 br_0_179 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c179
*+ bl_0_179 br_0_179 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c179
*+ bl_0_179 br_0_179 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c179
*+ bl_0_179 br_0_179 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c179
*+ bl_0_179 br_0_179 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c179
*+ bl_0_179 br_0_179 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c179
*+ bl_0_179 br_0_179 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c179
*+ bl_0_179 br_0_179 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c179
*+ bl_0_179 br_0_179 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c179
*+ bl_0_179 br_0_179 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c179
*+ bl_0_179 br_0_179 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c179
*+ bl_0_179 br_0_179 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c179
*+ bl_0_179 br_0_179 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c179
*+ bl_0_179 br_0_179 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c179
*+ bl_0_179 br_0_179 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c179
*+ bl_0_179 br_0_179 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c179
*+ bl_0_179 br_0_179 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c179
*+ bl_0_179 br_0_179 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c179
*+ bl_0_179 br_0_179 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c179
*+ bl_0_179 br_0_179 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c179
*+ bl_0_179 br_0_179 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c179
*+ bl_0_179 br_0_179 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c179
*+ bl_0_179 br_0_179 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c179
*+ bl_0_179 br_0_179 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c179
*+ bl_0_179 br_0_179 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c179
*+ bl_0_179 br_0_179 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c179
*+ bl_0_179 br_0_179 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c179
*+ bl_0_179 br_0_179 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c179
*+ bl_0_179 br_0_179 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c179
*+ bl_0_179 br_0_179 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c179
*+ bl_0_179 br_0_179 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c179
*+ bl_0_179 br_0_179 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c179
+ bl_0_179 br_0_179 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c180
+ bl_0_180 br_0_180 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c180
*+ bl_0_180 br_0_180 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c180
*+ bl_0_180 br_0_180 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c180
*+ bl_0_180 br_0_180 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c180
*+ bl_0_180 br_0_180 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c180
*+ bl_0_180 br_0_180 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c180
*+ bl_0_180 br_0_180 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c180
*+ bl_0_180 br_0_180 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c180
*+ bl_0_180 br_0_180 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c180
*+ bl_0_180 br_0_180 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c180
*+ bl_0_180 br_0_180 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c180
*+ bl_0_180 br_0_180 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c180
*+ bl_0_180 br_0_180 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c180
*+ bl_0_180 br_0_180 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c180
*+ bl_0_180 br_0_180 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c180
*+ bl_0_180 br_0_180 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c180
*+ bl_0_180 br_0_180 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c180
*+ bl_0_180 br_0_180 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c180
*+ bl_0_180 br_0_180 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c180
*+ bl_0_180 br_0_180 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c180
*+ bl_0_180 br_0_180 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c180
*+ bl_0_180 br_0_180 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c180
*+ bl_0_180 br_0_180 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c180
*+ bl_0_180 br_0_180 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c180
*+ bl_0_180 br_0_180 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c180
*+ bl_0_180 br_0_180 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c180
*+ bl_0_180 br_0_180 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c180
*+ bl_0_180 br_0_180 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c180
*+ bl_0_180 br_0_180 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c180
*+ bl_0_180 br_0_180 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c180
*+ bl_0_180 br_0_180 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c180
*+ bl_0_180 br_0_180 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c180
*+ bl_0_180 br_0_180 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c180
*+ bl_0_180 br_0_180 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c180
*+ bl_0_180 br_0_180 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c180
*+ bl_0_180 br_0_180 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c180
*+ bl_0_180 br_0_180 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c180
*+ bl_0_180 br_0_180 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c180
*+ bl_0_180 br_0_180 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c180
*+ bl_0_180 br_0_180 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c180
*+ bl_0_180 br_0_180 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c180
*+ bl_0_180 br_0_180 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c180
*+ bl_0_180 br_0_180 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c180
*+ bl_0_180 br_0_180 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c180
*+ bl_0_180 br_0_180 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c180
*+ bl_0_180 br_0_180 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c180
*+ bl_0_180 br_0_180 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c180
*+ bl_0_180 br_0_180 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c180
*+ bl_0_180 br_0_180 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c180
*+ bl_0_180 br_0_180 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c180
*+ bl_0_180 br_0_180 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c180
*+ bl_0_180 br_0_180 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c180
*+ bl_0_180 br_0_180 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c180
*+ bl_0_180 br_0_180 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c180
*+ bl_0_180 br_0_180 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c180
*+ bl_0_180 br_0_180 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c180
*+ bl_0_180 br_0_180 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c180
*+ bl_0_180 br_0_180 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c180
*+ bl_0_180 br_0_180 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c180
*+ bl_0_180 br_0_180 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c180
*+ bl_0_180 br_0_180 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c180
*+ bl_0_180 br_0_180 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c180
*+ bl_0_180 br_0_180 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c180
*+ bl_0_180 br_0_180 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c180
*+ bl_0_180 br_0_180 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c180
*+ bl_0_180 br_0_180 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c180
*+ bl_0_180 br_0_180 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c180
*+ bl_0_180 br_0_180 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c180
*+ bl_0_180 br_0_180 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c180
*+ bl_0_180 br_0_180 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c180
*+ bl_0_180 br_0_180 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c180
*+ bl_0_180 br_0_180 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c180
*+ bl_0_180 br_0_180 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c180
*+ bl_0_180 br_0_180 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c180
*+ bl_0_180 br_0_180 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c180
*+ bl_0_180 br_0_180 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c180
*+ bl_0_180 br_0_180 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c180
*+ bl_0_180 br_0_180 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c180
*+ bl_0_180 br_0_180 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c180
*+ bl_0_180 br_0_180 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c180
*+ bl_0_180 br_0_180 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c180
*+ bl_0_180 br_0_180 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c180
*+ bl_0_180 br_0_180 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c180
*+ bl_0_180 br_0_180 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c180
*+ bl_0_180 br_0_180 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c180
*+ bl_0_180 br_0_180 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c180
*+ bl_0_180 br_0_180 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c180
*+ bl_0_180 br_0_180 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c180
*+ bl_0_180 br_0_180 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c180
*+ bl_0_180 br_0_180 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c180
*+ bl_0_180 br_0_180 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c180
*+ bl_0_180 br_0_180 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c180
*+ bl_0_180 br_0_180 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c180
*+ bl_0_180 br_0_180 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c180
*+ bl_0_180 br_0_180 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c180
*+ bl_0_180 br_0_180 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c180
*+ bl_0_180 br_0_180 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c180
*+ bl_0_180 br_0_180 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c180
*+ bl_0_180 br_0_180 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c180
*+ bl_0_180 br_0_180 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c180
*+ bl_0_180 br_0_180 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c180
*+ bl_0_180 br_0_180 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c180
*+ bl_0_180 br_0_180 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c180
*+ bl_0_180 br_0_180 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c180
*+ bl_0_180 br_0_180 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c180
*+ bl_0_180 br_0_180 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c180
*+ bl_0_180 br_0_180 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c180
*+ bl_0_180 br_0_180 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c180
*+ bl_0_180 br_0_180 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c180
*+ bl_0_180 br_0_180 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c180
*+ bl_0_180 br_0_180 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c180
*+ bl_0_180 br_0_180 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c180
*+ bl_0_180 br_0_180 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c180
*+ bl_0_180 br_0_180 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c180
*+ bl_0_180 br_0_180 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c180
*+ bl_0_180 br_0_180 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c180
*+ bl_0_180 br_0_180 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c180
*+ bl_0_180 br_0_180 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c180
*+ bl_0_180 br_0_180 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c180
*+ bl_0_180 br_0_180 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c180
*+ bl_0_180 br_0_180 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c180
*+ bl_0_180 br_0_180 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c180
*+ bl_0_180 br_0_180 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c180
*+ bl_0_180 br_0_180 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c180
*+ bl_0_180 br_0_180 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c180
*+ bl_0_180 br_0_180 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c180
*+ bl_0_180 br_0_180 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c180
+ bl_0_180 br_0_180 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c181
+ bl_0_181 br_0_181 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c181
*+ bl_0_181 br_0_181 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c181
*+ bl_0_181 br_0_181 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c181
*+ bl_0_181 br_0_181 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c181
*+ bl_0_181 br_0_181 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c181
*+ bl_0_181 br_0_181 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c181
*+ bl_0_181 br_0_181 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c181
*+ bl_0_181 br_0_181 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c181
*+ bl_0_181 br_0_181 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c181
*+ bl_0_181 br_0_181 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c181
*+ bl_0_181 br_0_181 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c181
*+ bl_0_181 br_0_181 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c181
*+ bl_0_181 br_0_181 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c181
*+ bl_0_181 br_0_181 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c181
*+ bl_0_181 br_0_181 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c181
*+ bl_0_181 br_0_181 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c181
*+ bl_0_181 br_0_181 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c181
*+ bl_0_181 br_0_181 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c181
*+ bl_0_181 br_0_181 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c181
*+ bl_0_181 br_0_181 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c181
*+ bl_0_181 br_0_181 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c181
*+ bl_0_181 br_0_181 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c181
*+ bl_0_181 br_0_181 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c181
*+ bl_0_181 br_0_181 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c181
*+ bl_0_181 br_0_181 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c181
*+ bl_0_181 br_0_181 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c181
*+ bl_0_181 br_0_181 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c181
*+ bl_0_181 br_0_181 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c181
*+ bl_0_181 br_0_181 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c181
*+ bl_0_181 br_0_181 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c181
*+ bl_0_181 br_0_181 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c181
*+ bl_0_181 br_0_181 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c181
*+ bl_0_181 br_0_181 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c181
*+ bl_0_181 br_0_181 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c181
*+ bl_0_181 br_0_181 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c181
*+ bl_0_181 br_0_181 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c181
*+ bl_0_181 br_0_181 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c181
*+ bl_0_181 br_0_181 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c181
*+ bl_0_181 br_0_181 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c181
*+ bl_0_181 br_0_181 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c181
*+ bl_0_181 br_0_181 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c181
*+ bl_0_181 br_0_181 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c181
*+ bl_0_181 br_0_181 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c181
*+ bl_0_181 br_0_181 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c181
*+ bl_0_181 br_0_181 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c181
*+ bl_0_181 br_0_181 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c181
*+ bl_0_181 br_0_181 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c181
*+ bl_0_181 br_0_181 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c181
*+ bl_0_181 br_0_181 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c181
*+ bl_0_181 br_0_181 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c181
*+ bl_0_181 br_0_181 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c181
*+ bl_0_181 br_0_181 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c181
*+ bl_0_181 br_0_181 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c181
*+ bl_0_181 br_0_181 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c181
*+ bl_0_181 br_0_181 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c181
*+ bl_0_181 br_0_181 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c181
*+ bl_0_181 br_0_181 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c181
*+ bl_0_181 br_0_181 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c181
*+ bl_0_181 br_0_181 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c181
*+ bl_0_181 br_0_181 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c181
*+ bl_0_181 br_0_181 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c181
*+ bl_0_181 br_0_181 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c181
*+ bl_0_181 br_0_181 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c181
*+ bl_0_181 br_0_181 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c181
*+ bl_0_181 br_0_181 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c181
*+ bl_0_181 br_0_181 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c181
*+ bl_0_181 br_0_181 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c181
*+ bl_0_181 br_0_181 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c181
*+ bl_0_181 br_0_181 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c181
*+ bl_0_181 br_0_181 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c181
*+ bl_0_181 br_0_181 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c181
*+ bl_0_181 br_0_181 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c181
*+ bl_0_181 br_0_181 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c181
*+ bl_0_181 br_0_181 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c181
*+ bl_0_181 br_0_181 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c181
*+ bl_0_181 br_0_181 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c181
*+ bl_0_181 br_0_181 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c181
*+ bl_0_181 br_0_181 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c181
*+ bl_0_181 br_0_181 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c181
*+ bl_0_181 br_0_181 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c181
*+ bl_0_181 br_0_181 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c181
*+ bl_0_181 br_0_181 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c181
*+ bl_0_181 br_0_181 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c181
*+ bl_0_181 br_0_181 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c181
*+ bl_0_181 br_0_181 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c181
*+ bl_0_181 br_0_181 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c181
*+ bl_0_181 br_0_181 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c181
*+ bl_0_181 br_0_181 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c181
*+ bl_0_181 br_0_181 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c181
*+ bl_0_181 br_0_181 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c181
*+ bl_0_181 br_0_181 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c181
*+ bl_0_181 br_0_181 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c181
*+ bl_0_181 br_0_181 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c181
*+ bl_0_181 br_0_181 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c181
*+ bl_0_181 br_0_181 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c181
*+ bl_0_181 br_0_181 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c181
*+ bl_0_181 br_0_181 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c181
*+ bl_0_181 br_0_181 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c181
*+ bl_0_181 br_0_181 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c181
*+ bl_0_181 br_0_181 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c181
*+ bl_0_181 br_0_181 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c181
*+ bl_0_181 br_0_181 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c181
*+ bl_0_181 br_0_181 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c181
*+ bl_0_181 br_0_181 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c181
*+ bl_0_181 br_0_181 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c181
*+ bl_0_181 br_0_181 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c181
*+ bl_0_181 br_0_181 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c181
*+ bl_0_181 br_0_181 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c181
*+ bl_0_181 br_0_181 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c181
*+ bl_0_181 br_0_181 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c181
*+ bl_0_181 br_0_181 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c181
*+ bl_0_181 br_0_181 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c181
*+ bl_0_181 br_0_181 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c181
*+ bl_0_181 br_0_181 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c181
*+ bl_0_181 br_0_181 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c181
*+ bl_0_181 br_0_181 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c181
*+ bl_0_181 br_0_181 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c181
*+ bl_0_181 br_0_181 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c181
*+ bl_0_181 br_0_181 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c181
*+ bl_0_181 br_0_181 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c181
*+ bl_0_181 br_0_181 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c181
*+ bl_0_181 br_0_181 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c181
*+ bl_0_181 br_0_181 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c181
*+ bl_0_181 br_0_181 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c181
*+ bl_0_181 br_0_181 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c181
*+ bl_0_181 br_0_181 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c181
*+ bl_0_181 br_0_181 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c181
+ bl_0_181 br_0_181 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c182
+ bl_0_182 br_0_182 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c182
*+ bl_0_182 br_0_182 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c182
*+ bl_0_182 br_0_182 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c182
*+ bl_0_182 br_0_182 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c182
*+ bl_0_182 br_0_182 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c182
*+ bl_0_182 br_0_182 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c182
*+ bl_0_182 br_0_182 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c182
*+ bl_0_182 br_0_182 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c182
*+ bl_0_182 br_0_182 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c182
*+ bl_0_182 br_0_182 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c182
*+ bl_0_182 br_0_182 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c182
*+ bl_0_182 br_0_182 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c182
*+ bl_0_182 br_0_182 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c182
*+ bl_0_182 br_0_182 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c182
*+ bl_0_182 br_0_182 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c182
*+ bl_0_182 br_0_182 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c182
*+ bl_0_182 br_0_182 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c182
*+ bl_0_182 br_0_182 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c182
*+ bl_0_182 br_0_182 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c182
*+ bl_0_182 br_0_182 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c182
*+ bl_0_182 br_0_182 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c182
*+ bl_0_182 br_0_182 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c182
*+ bl_0_182 br_0_182 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c182
*+ bl_0_182 br_0_182 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c182
*+ bl_0_182 br_0_182 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c182
*+ bl_0_182 br_0_182 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c182
*+ bl_0_182 br_0_182 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c182
*+ bl_0_182 br_0_182 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c182
*+ bl_0_182 br_0_182 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c182
*+ bl_0_182 br_0_182 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c182
*+ bl_0_182 br_0_182 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c182
*+ bl_0_182 br_0_182 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c182
*+ bl_0_182 br_0_182 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c182
*+ bl_0_182 br_0_182 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c182
*+ bl_0_182 br_0_182 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c182
*+ bl_0_182 br_0_182 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c182
*+ bl_0_182 br_0_182 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c182
*+ bl_0_182 br_0_182 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c182
*+ bl_0_182 br_0_182 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c182
*+ bl_0_182 br_0_182 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c182
*+ bl_0_182 br_0_182 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c182
*+ bl_0_182 br_0_182 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c182
*+ bl_0_182 br_0_182 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c182
*+ bl_0_182 br_0_182 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c182
*+ bl_0_182 br_0_182 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c182
*+ bl_0_182 br_0_182 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c182
*+ bl_0_182 br_0_182 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c182
*+ bl_0_182 br_0_182 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c182
*+ bl_0_182 br_0_182 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c182
*+ bl_0_182 br_0_182 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c182
*+ bl_0_182 br_0_182 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c182
*+ bl_0_182 br_0_182 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c182
*+ bl_0_182 br_0_182 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c182
*+ bl_0_182 br_0_182 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c182
*+ bl_0_182 br_0_182 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c182
*+ bl_0_182 br_0_182 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c182
*+ bl_0_182 br_0_182 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c182
*+ bl_0_182 br_0_182 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c182
*+ bl_0_182 br_0_182 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c182
*+ bl_0_182 br_0_182 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c182
*+ bl_0_182 br_0_182 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c182
*+ bl_0_182 br_0_182 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c182
*+ bl_0_182 br_0_182 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c182
*+ bl_0_182 br_0_182 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c182
*+ bl_0_182 br_0_182 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c182
*+ bl_0_182 br_0_182 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c182
*+ bl_0_182 br_0_182 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c182
*+ bl_0_182 br_0_182 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c182
*+ bl_0_182 br_0_182 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c182
*+ bl_0_182 br_0_182 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c182
*+ bl_0_182 br_0_182 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c182
*+ bl_0_182 br_0_182 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c182
*+ bl_0_182 br_0_182 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c182
*+ bl_0_182 br_0_182 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c182
*+ bl_0_182 br_0_182 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c182
*+ bl_0_182 br_0_182 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c182
*+ bl_0_182 br_0_182 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c182
*+ bl_0_182 br_0_182 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c182
*+ bl_0_182 br_0_182 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c182
*+ bl_0_182 br_0_182 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c182
*+ bl_0_182 br_0_182 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c182
*+ bl_0_182 br_0_182 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c182
*+ bl_0_182 br_0_182 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c182
*+ bl_0_182 br_0_182 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c182
*+ bl_0_182 br_0_182 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c182
*+ bl_0_182 br_0_182 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c182
*+ bl_0_182 br_0_182 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c182
*+ bl_0_182 br_0_182 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c182
*+ bl_0_182 br_0_182 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c182
*+ bl_0_182 br_0_182 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c182
*+ bl_0_182 br_0_182 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c182
*+ bl_0_182 br_0_182 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c182
*+ bl_0_182 br_0_182 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c182
*+ bl_0_182 br_0_182 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c182
*+ bl_0_182 br_0_182 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c182
*+ bl_0_182 br_0_182 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c182
*+ bl_0_182 br_0_182 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c182
*+ bl_0_182 br_0_182 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c182
*+ bl_0_182 br_0_182 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c182
*+ bl_0_182 br_0_182 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c182
*+ bl_0_182 br_0_182 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c182
*+ bl_0_182 br_0_182 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c182
*+ bl_0_182 br_0_182 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c182
*+ bl_0_182 br_0_182 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c182
*+ bl_0_182 br_0_182 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c182
*+ bl_0_182 br_0_182 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c182
*+ bl_0_182 br_0_182 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c182
*+ bl_0_182 br_0_182 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c182
*+ bl_0_182 br_0_182 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c182
*+ bl_0_182 br_0_182 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c182
*+ bl_0_182 br_0_182 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c182
*+ bl_0_182 br_0_182 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c182
*+ bl_0_182 br_0_182 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c182
*+ bl_0_182 br_0_182 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c182
*+ bl_0_182 br_0_182 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c182
*+ bl_0_182 br_0_182 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c182
*+ bl_0_182 br_0_182 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c182
*+ bl_0_182 br_0_182 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c182
*+ bl_0_182 br_0_182 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c182
*+ bl_0_182 br_0_182 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c182
*+ bl_0_182 br_0_182 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c182
*+ bl_0_182 br_0_182 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c182
*+ bl_0_182 br_0_182 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c182
*+ bl_0_182 br_0_182 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c182
*+ bl_0_182 br_0_182 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c182
*+ bl_0_182 br_0_182 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c182
*+ bl_0_182 br_0_182 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c182
+ bl_0_182 br_0_182 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c183
+ bl_0_183 br_0_183 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c183
*+ bl_0_183 br_0_183 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c183
*+ bl_0_183 br_0_183 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c183
*+ bl_0_183 br_0_183 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c183
*+ bl_0_183 br_0_183 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c183
*+ bl_0_183 br_0_183 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c183
*+ bl_0_183 br_0_183 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c183
*+ bl_0_183 br_0_183 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c183
*+ bl_0_183 br_0_183 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c183
*+ bl_0_183 br_0_183 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c183
*+ bl_0_183 br_0_183 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c183
*+ bl_0_183 br_0_183 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c183
*+ bl_0_183 br_0_183 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c183
*+ bl_0_183 br_0_183 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c183
*+ bl_0_183 br_0_183 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c183
*+ bl_0_183 br_0_183 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c183
*+ bl_0_183 br_0_183 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c183
*+ bl_0_183 br_0_183 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c183
*+ bl_0_183 br_0_183 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c183
*+ bl_0_183 br_0_183 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c183
*+ bl_0_183 br_0_183 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c183
*+ bl_0_183 br_0_183 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c183
*+ bl_0_183 br_0_183 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c183
*+ bl_0_183 br_0_183 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c183
*+ bl_0_183 br_0_183 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c183
*+ bl_0_183 br_0_183 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c183
*+ bl_0_183 br_0_183 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c183
*+ bl_0_183 br_0_183 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c183
*+ bl_0_183 br_0_183 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c183
*+ bl_0_183 br_0_183 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c183
*+ bl_0_183 br_0_183 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c183
*+ bl_0_183 br_0_183 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c183
*+ bl_0_183 br_0_183 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c183
*+ bl_0_183 br_0_183 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c183
*+ bl_0_183 br_0_183 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c183
*+ bl_0_183 br_0_183 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c183
*+ bl_0_183 br_0_183 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c183
*+ bl_0_183 br_0_183 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c183
*+ bl_0_183 br_0_183 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c183
*+ bl_0_183 br_0_183 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c183
*+ bl_0_183 br_0_183 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c183
*+ bl_0_183 br_0_183 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c183
*+ bl_0_183 br_0_183 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c183
*+ bl_0_183 br_0_183 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c183
*+ bl_0_183 br_0_183 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c183
*+ bl_0_183 br_0_183 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c183
*+ bl_0_183 br_0_183 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c183
*+ bl_0_183 br_0_183 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c183
*+ bl_0_183 br_0_183 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c183
*+ bl_0_183 br_0_183 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c183
*+ bl_0_183 br_0_183 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c183
*+ bl_0_183 br_0_183 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c183
*+ bl_0_183 br_0_183 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c183
*+ bl_0_183 br_0_183 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c183
*+ bl_0_183 br_0_183 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c183
*+ bl_0_183 br_0_183 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c183
*+ bl_0_183 br_0_183 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c183
*+ bl_0_183 br_0_183 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c183
*+ bl_0_183 br_0_183 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c183
*+ bl_0_183 br_0_183 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c183
*+ bl_0_183 br_0_183 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c183
*+ bl_0_183 br_0_183 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c183
*+ bl_0_183 br_0_183 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c183
*+ bl_0_183 br_0_183 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c183
*+ bl_0_183 br_0_183 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c183
*+ bl_0_183 br_0_183 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c183
*+ bl_0_183 br_0_183 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c183
*+ bl_0_183 br_0_183 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c183
*+ bl_0_183 br_0_183 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c183
*+ bl_0_183 br_0_183 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c183
*+ bl_0_183 br_0_183 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c183
*+ bl_0_183 br_0_183 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c183
*+ bl_0_183 br_0_183 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c183
*+ bl_0_183 br_0_183 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c183
*+ bl_0_183 br_0_183 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c183
*+ bl_0_183 br_0_183 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c183
*+ bl_0_183 br_0_183 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c183
*+ bl_0_183 br_0_183 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c183
*+ bl_0_183 br_0_183 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c183
*+ bl_0_183 br_0_183 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c183
*+ bl_0_183 br_0_183 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c183
*+ bl_0_183 br_0_183 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c183
*+ bl_0_183 br_0_183 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c183
*+ bl_0_183 br_0_183 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c183
*+ bl_0_183 br_0_183 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c183
*+ bl_0_183 br_0_183 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c183
*+ bl_0_183 br_0_183 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c183
*+ bl_0_183 br_0_183 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c183
*+ bl_0_183 br_0_183 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c183
*+ bl_0_183 br_0_183 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c183
*+ bl_0_183 br_0_183 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c183
*+ bl_0_183 br_0_183 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c183
*+ bl_0_183 br_0_183 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c183
*+ bl_0_183 br_0_183 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c183
*+ bl_0_183 br_0_183 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c183
*+ bl_0_183 br_0_183 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c183
*+ bl_0_183 br_0_183 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c183
*+ bl_0_183 br_0_183 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c183
*+ bl_0_183 br_0_183 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c183
*+ bl_0_183 br_0_183 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c183
*+ bl_0_183 br_0_183 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c183
*+ bl_0_183 br_0_183 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c183
*+ bl_0_183 br_0_183 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c183
*+ bl_0_183 br_0_183 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c183
*+ bl_0_183 br_0_183 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c183
*+ bl_0_183 br_0_183 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c183
*+ bl_0_183 br_0_183 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c183
*+ bl_0_183 br_0_183 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c183
*+ bl_0_183 br_0_183 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c183
*+ bl_0_183 br_0_183 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c183
*+ bl_0_183 br_0_183 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c183
*+ bl_0_183 br_0_183 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c183
*+ bl_0_183 br_0_183 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c183
*+ bl_0_183 br_0_183 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c183
*+ bl_0_183 br_0_183 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c183
*+ bl_0_183 br_0_183 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c183
*+ bl_0_183 br_0_183 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c183
*+ bl_0_183 br_0_183 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c183
*+ bl_0_183 br_0_183 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c183
*+ bl_0_183 br_0_183 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c183
*+ bl_0_183 br_0_183 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c183
*+ bl_0_183 br_0_183 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c183
*+ bl_0_183 br_0_183 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c183
*+ bl_0_183 br_0_183 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c183
*+ bl_0_183 br_0_183 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c183
*+ bl_0_183 br_0_183 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c183
*+ bl_0_183 br_0_183 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c183
+ bl_0_183 br_0_183 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c184
+ bl_0_184 br_0_184 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c184
*+ bl_0_184 br_0_184 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c184
*+ bl_0_184 br_0_184 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c184
*+ bl_0_184 br_0_184 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c184
*+ bl_0_184 br_0_184 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c184
*+ bl_0_184 br_0_184 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c184
*+ bl_0_184 br_0_184 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c184
*+ bl_0_184 br_0_184 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c184
*+ bl_0_184 br_0_184 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c184
*+ bl_0_184 br_0_184 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c184
*+ bl_0_184 br_0_184 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c184
*+ bl_0_184 br_0_184 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c184
*+ bl_0_184 br_0_184 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c184
*+ bl_0_184 br_0_184 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c184
*+ bl_0_184 br_0_184 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c184
*+ bl_0_184 br_0_184 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c184
*+ bl_0_184 br_0_184 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c184
*+ bl_0_184 br_0_184 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c184
*+ bl_0_184 br_0_184 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c184
*+ bl_0_184 br_0_184 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c184
*+ bl_0_184 br_0_184 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c184
*+ bl_0_184 br_0_184 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c184
*+ bl_0_184 br_0_184 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c184
*+ bl_0_184 br_0_184 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c184
*+ bl_0_184 br_0_184 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c184
*+ bl_0_184 br_0_184 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c184
*+ bl_0_184 br_0_184 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c184
*+ bl_0_184 br_0_184 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c184
*+ bl_0_184 br_0_184 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c184
*+ bl_0_184 br_0_184 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c184
*+ bl_0_184 br_0_184 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c184
*+ bl_0_184 br_0_184 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c184
*+ bl_0_184 br_0_184 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c184
*+ bl_0_184 br_0_184 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c184
*+ bl_0_184 br_0_184 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c184
*+ bl_0_184 br_0_184 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c184
*+ bl_0_184 br_0_184 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c184
*+ bl_0_184 br_0_184 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c184
*+ bl_0_184 br_0_184 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c184
*+ bl_0_184 br_0_184 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c184
*+ bl_0_184 br_0_184 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c184
*+ bl_0_184 br_0_184 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c184
*+ bl_0_184 br_0_184 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c184
*+ bl_0_184 br_0_184 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c184
*+ bl_0_184 br_0_184 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c184
*+ bl_0_184 br_0_184 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c184
*+ bl_0_184 br_0_184 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c184
*+ bl_0_184 br_0_184 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c184
*+ bl_0_184 br_0_184 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c184
*+ bl_0_184 br_0_184 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c184
*+ bl_0_184 br_0_184 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c184
*+ bl_0_184 br_0_184 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c184
*+ bl_0_184 br_0_184 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c184
*+ bl_0_184 br_0_184 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c184
*+ bl_0_184 br_0_184 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c184
*+ bl_0_184 br_0_184 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c184
*+ bl_0_184 br_0_184 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c184
*+ bl_0_184 br_0_184 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c184
*+ bl_0_184 br_0_184 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c184
*+ bl_0_184 br_0_184 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c184
*+ bl_0_184 br_0_184 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c184
*+ bl_0_184 br_0_184 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c184
*+ bl_0_184 br_0_184 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c184
*+ bl_0_184 br_0_184 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c184
*+ bl_0_184 br_0_184 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c184
*+ bl_0_184 br_0_184 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c184
*+ bl_0_184 br_0_184 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c184
*+ bl_0_184 br_0_184 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c184
*+ bl_0_184 br_0_184 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c184
*+ bl_0_184 br_0_184 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c184
*+ bl_0_184 br_0_184 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c184
*+ bl_0_184 br_0_184 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c184
*+ bl_0_184 br_0_184 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c184
*+ bl_0_184 br_0_184 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c184
*+ bl_0_184 br_0_184 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c184
*+ bl_0_184 br_0_184 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c184
*+ bl_0_184 br_0_184 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c184
*+ bl_0_184 br_0_184 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c184
*+ bl_0_184 br_0_184 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c184
*+ bl_0_184 br_0_184 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c184
*+ bl_0_184 br_0_184 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c184
*+ bl_0_184 br_0_184 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c184
*+ bl_0_184 br_0_184 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c184
*+ bl_0_184 br_0_184 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c184
*+ bl_0_184 br_0_184 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c184
*+ bl_0_184 br_0_184 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c184
*+ bl_0_184 br_0_184 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c184
*+ bl_0_184 br_0_184 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c184
*+ bl_0_184 br_0_184 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c184
*+ bl_0_184 br_0_184 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c184
*+ bl_0_184 br_0_184 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c184
*+ bl_0_184 br_0_184 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c184
*+ bl_0_184 br_0_184 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c184
*+ bl_0_184 br_0_184 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c184
*+ bl_0_184 br_0_184 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c184
*+ bl_0_184 br_0_184 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c184
*+ bl_0_184 br_0_184 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c184
*+ bl_0_184 br_0_184 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c184
*+ bl_0_184 br_0_184 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c184
*+ bl_0_184 br_0_184 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c184
*+ bl_0_184 br_0_184 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c184
*+ bl_0_184 br_0_184 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c184
*+ bl_0_184 br_0_184 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c184
*+ bl_0_184 br_0_184 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c184
*+ bl_0_184 br_0_184 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c184
*+ bl_0_184 br_0_184 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c184
*+ bl_0_184 br_0_184 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c184
*+ bl_0_184 br_0_184 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c184
*+ bl_0_184 br_0_184 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c184
*+ bl_0_184 br_0_184 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c184
*+ bl_0_184 br_0_184 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c184
*+ bl_0_184 br_0_184 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c184
*+ bl_0_184 br_0_184 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c184
*+ bl_0_184 br_0_184 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c184
*+ bl_0_184 br_0_184 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c184
*+ bl_0_184 br_0_184 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c184
*+ bl_0_184 br_0_184 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c184
*+ bl_0_184 br_0_184 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c184
*+ bl_0_184 br_0_184 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c184
*+ bl_0_184 br_0_184 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c184
*+ bl_0_184 br_0_184 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c184
*+ bl_0_184 br_0_184 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c184
*+ bl_0_184 br_0_184 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c184
*+ bl_0_184 br_0_184 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c184
*+ bl_0_184 br_0_184 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c184
*+ bl_0_184 br_0_184 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c184
*+ bl_0_184 br_0_184 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c184
+ bl_0_184 br_0_184 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c185
+ bl_0_185 br_0_185 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c185
*+ bl_0_185 br_0_185 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c185
*+ bl_0_185 br_0_185 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c185
*+ bl_0_185 br_0_185 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c185
*+ bl_0_185 br_0_185 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c185
*+ bl_0_185 br_0_185 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c185
*+ bl_0_185 br_0_185 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c185
*+ bl_0_185 br_0_185 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c185
*+ bl_0_185 br_0_185 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c185
*+ bl_0_185 br_0_185 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c185
*+ bl_0_185 br_0_185 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c185
*+ bl_0_185 br_0_185 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c185
*+ bl_0_185 br_0_185 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c185
*+ bl_0_185 br_0_185 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c185
*+ bl_0_185 br_0_185 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c185
*+ bl_0_185 br_0_185 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c185
*+ bl_0_185 br_0_185 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c185
*+ bl_0_185 br_0_185 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c185
*+ bl_0_185 br_0_185 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c185
*+ bl_0_185 br_0_185 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c185
*+ bl_0_185 br_0_185 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c185
*+ bl_0_185 br_0_185 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c185
*+ bl_0_185 br_0_185 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c185
*+ bl_0_185 br_0_185 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c185
*+ bl_0_185 br_0_185 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c185
*+ bl_0_185 br_0_185 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c185
*+ bl_0_185 br_0_185 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c185
*+ bl_0_185 br_0_185 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c185
*+ bl_0_185 br_0_185 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c185
*+ bl_0_185 br_0_185 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c185
*+ bl_0_185 br_0_185 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c185
*+ bl_0_185 br_0_185 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c185
*+ bl_0_185 br_0_185 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c185
*+ bl_0_185 br_0_185 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c185
*+ bl_0_185 br_0_185 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c185
*+ bl_0_185 br_0_185 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c185
*+ bl_0_185 br_0_185 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c185
*+ bl_0_185 br_0_185 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c185
*+ bl_0_185 br_0_185 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c185
*+ bl_0_185 br_0_185 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c185
*+ bl_0_185 br_0_185 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c185
*+ bl_0_185 br_0_185 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c185
*+ bl_0_185 br_0_185 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c185
*+ bl_0_185 br_0_185 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c185
*+ bl_0_185 br_0_185 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c185
*+ bl_0_185 br_0_185 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c185
*+ bl_0_185 br_0_185 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c185
*+ bl_0_185 br_0_185 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c185
*+ bl_0_185 br_0_185 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c185
*+ bl_0_185 br_0_185 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c185
*+ bl_0_185 br_0_185 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c185
*+ bl_0_185 br_0_185 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c185
*+ bl_0_185 br_0_185 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c185
*+ bl_0_185 br_0_185 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c185
*+ bl_0_185 br_0_185 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c185
*+ bl_0_185 br_0_185 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c185
*+ bl_0_185 br_0_185 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c185
*+ bl_0_185 br_0_185 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c185
*+ bl_0_185 br_0_185 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c185
*+ bl_0_185 br_0_185 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c185
*+ bl_0_185 br_0_185 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c185
*+ bl_0_185 br_0_185 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c185
*+ bl_0_185 br_0_185 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c185
*+ bl_0_185 br_0_185 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c185
*+ bl_0_185 br_0_185 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c185
*+ bl_0_185 br_0_185 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c185
*+ bl_0_185 br_0_185 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c185
*+ bl_0_185 br_0_185 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c185
*+ bl_0_185 br_0_185 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c185
*+ bl_0_185 br_0_185 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c185
*+ bl_0_185 br_0_185 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c185
*+ bl_0_185 br_0_185 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c185
*+ bl_0_185 br_0_185 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c185
*+ bl_0_185 br_0_185 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c185
*+ bl_0_185 br_0_185 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c185
*+ bl_0_185 br_0_185 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c185
*+ bl_0_185 br_0_185 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c185
*+ bl_0_185 br_0_185 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c185
*+ bl_0_185 br_0_185 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c185
*+ bl_0_185 br_0_185 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c185
*+ bl_0_185 br_0_185 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c185
*+ bl_0_185 br_0_185 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c185
*+ bl_0_185 br_0_185 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c185
*+ bl_0_185 br_0_185 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c185
*+ bl_0_185 br_0_185 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c185
*+ bl_0_185 br_0_185 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c185
*+ bl_0_185 br_0_185 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c185
*+ bl_0_185 br_0_185 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c185
*+ bl_0_185 br_0_185 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c185
*+ bl_0_185 br_0_185 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c185
*+ bl_0_185 br_0_185 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c185
*+ bl_0_185 br_0_185 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c185
*+ bl_0_185 br_0_185 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c185
*+ bl_0_185 br_0_185 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c185
*+ bl_0_185 br_0_185 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c185
*+ bl_0_185 br_0_185 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c185
*+ bl_0_185 br_0_185 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c185
*+ bl_0_185 br_0_185 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c185
*+ bl_0_185 br_0_185 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c185
*+ bl_0_185 br_0_185 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c185
*+ bl_0_185 br_0_185 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c185
*+ bl_0_185 br_0_185 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c185
*+ bl_0_185 br_0_185 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c185
*+ bl_0_185 br_0_185 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c185
*+ bl_0_185 br_0_185 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c185
*+ bl_0_185 br_0_185 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c185
*+ bl_0_185 br_0_185 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c185
*+ bl_0_185 br_0_185 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c185
*+ bl_0_185 br_0_185 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c185
*+ bl_0_185 br_0_185 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c185
*+ bl_0_185 br_0_185 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c185
*+ bl_0_185 br_0_185 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c185
*+ bl_0_185 br_0_185 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c185
*+ bl_0_185 br_0_185 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c185
*+ bl_0_185 br_0_185 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c185
*+ bl_0_185 br_0_185 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c185
*+ bl_0_185 br_0_185 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c185
*+ bl_0_185 br_0_185 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c185
*+ bl_0_185 br_0_185 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c185
*+ bl_0_185 br_0_185 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c185
*+ bl_0_185 br_0_185 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c185
*+ bl_0_185 br_0_185 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c185
*+ bl_0_185 br_0_185 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c185
*+ bl_0_185 br_0_185 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c185
*+ bl_0_185 br_0_185 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c185
*+ bl_0_185 br_0_185 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c185
*+ bl_0_185 br_0_185 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c185
+ bl_0_185 br_0_185 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c186
+ bl_0_186 br_0_186 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c186
*+ bl_0_186 br_0_186 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c186
*+ bl_0_186 br_0_186 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c186
*+ bl_0_186 br_0_186 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c186
*+ bl_0_186 br_0_186 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c186
*+ bl_0_186 br_0_186 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c186
*+ bl_0_186 br_0_186 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c186
*+ bl_0_186 br_0_186 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c186
*+ bl_0_186 br_0_186 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c186
*+ bl_0_186 br_0_186 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c186
*+ bl_0_186 br_0_186 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c186
*+ bl_0_186 br_0_186 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c186
*+ bl_0_186 br_0_186 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c186
*+ bl_0_186 br_0_186 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c186
*+ bl_0_186 br_0_186 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c186
*+ bl_0_186 br_0_186 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c186
*+ bl_0_186 br_0_186 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c186
*+ bl_0_186 br_0_186 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c186
*+ bl_0_186 br_0_186 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c186
*+ bl_0_186 br_0_186 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c186
*+ bl_0_186 br_0_186 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c186
*+ bl_0_186 br_0_186 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c186
*+ bl_0_186 br_0_186 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c186
*+ bl_0_186 br_0_186 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c186
*+ bl_0_186 br_0_186 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c186
*+ bl_0_186 br_0_186 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c186
*+ bl_0_186 br_0_186 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c186
*+ bl_0_186 br_0_186 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c186
*+ bl_0_186 br_0_186 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c186
*+ bl_0_186 br_0_186 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c186
*+ bl_0_186 br_0_186 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c186
*+ bl_0_186 br_0_186 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c186
*+ bl_0_186 br_0_186 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c186
*+ bl_0_186 br_0_186 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c186
*+ bl_0_186 br_0_186 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c186
*+ bl_0_186 br_0_186 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c186
*+ bl_0_186 br_0_186 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c186
*+ bl_0_186 br_0_186 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c186
*+ bl_0_186 br_0_186 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c186
*+ bl_0_186 br_0_186 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c186
*+ bl_0_186 br_0_186 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c186
*+ bl_0_186 br_0_186 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c186
*+ bl_0_186 br_0_186 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c186
*+ bl_0_186 br_0_186 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c186
*+ bl_0_186 br_0_186 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c186
*+ bl_0_186 br_0_186 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c186
*+ bl_0_186 br_0_186 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c186
*+ bl_0_186 br_0_186 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c186
*+ bl_0_186 br_0_186 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c186
*+ bl_0_186 br_0_186 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c186
*+ bl_0_186 br_0_186 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c186
*+ bl_0_186 br_0_186 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c186
*+ bl_0_186 br_0_186 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c186
*+ bl_0_186 br_0_186 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c186
*+ bl_0_186 br_0_186 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c186
*+ bl_0_186 br_0_186 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c186
*+ bl_0_186 br_0_186 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c186
*+ bl_0_186 br_0_186 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c186
*+ bl_0_186 br_0_186 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c186
*+ bl_0_186 br_0_186 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c186
*+ bl_0_186 br_0_186 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c186
*+ bl_0_186 br_0_186 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c186
*+ bl_0_186 br_0_186 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c186
*+ bl_0_186 br_0_186 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c186
*+ bl_0_186 br_0_186 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c186
*+ bl_0_186 br_0_186 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c186
*+ bl_0_186 br_0_186 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c186
*+ bl_0_186 br_0_186 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c186
*+ bl_0_186 br_0_186 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c186
*+ bl_0_186 br_0_186 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c186
*+ bl_0_186 br_0_186 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c186
*+ bl_0_186 br_0_186 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c186
*+ bl_0_186 br_0_186 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c186
*+ bl_0_186 br_0_186 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c186
*+ bl_0_186 br_0_186 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c186
*+ bl_0_186 br_0_186 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c186
*+ bl_0_186 br_0_186 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c186
*+ bl_0_186 br_0_186 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c186
*+ bl_0_186 br_0_186 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c186
*+ bl_0_186 br_0_186 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c186
*+ bl_0_186 br_0_186 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c186
*+ bl_0_186 br_0_186 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c186
*+ bl_0_186 br_0_186 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c186
*+ bl_0_186 br_0_186 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c186
*+ bl_0_186 br_0_186 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c186
*+ bl_0_186 br_0_186 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c186
*+ bl_0_186 br_0_186 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c186
*+ bl_0_186 br_0_186 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c186
*+ bl_0_186 br_0_186 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c186
*+ bl_0_186 br_0_186 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c186
*+ bl_0_186 br_0_186 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c186
*+ bl_0_186 br_0_186 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c186
*+ bl_0_186 br_0_186 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c186
*+ bl_0_186 br_0_186 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c186
*+ bl_0_186 br_0_186 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c186
*+ bl_0_186 br_0_186 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c186
*+ bl_0_186 br_0_186 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c186
*+ bl_0_186 br_0_186 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c186
*+ bl_0_186 br_0_186 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c186
*+ bl_0_186 br_0_186 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c186
*+ bl_0_186 br_0_186 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c186
*+ bl_0_186 br_0_186 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c186
*+ bl_0_186 br_0_186 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c186
*+ bl_0_186 br_0_186 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c186
*+ bl_0_186 br_0_186 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c186
*+ bl_0_186 br_0_186 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c186
*+ bl_0_186 br_0_186 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c186
*+ bl_0_186 br_0_186 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c186
*+ bl_0_186 br_0_186 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c186
*+ bl_0_186 br_0_186 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c186
*+ bl_0_186 br_0_186 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c186
*+ bl_0_186 br_0_186 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c186
*+ bl_0_186 br_0_186 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c186
*+ bl_0_186 br_0_186 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c186
*+ bl_0_186 br_0_186 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c186
*+ bl_0_186 br_0_186 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c186
*+ bl_0_186 br_0_186 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c186
*+ bl_0_186 br_0_186 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c186
*+ bl_0_186 br_0_186 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c186
*+ bl_0_186 br_0_186 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c186
*+ bl_0_186 br_0_186 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c186
*+ bl_0_186 br_0_186 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c186
*+ bl_0_186 br_0_186 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c186
*+ bl_0_186 br_0_186 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c186
*+ bl_0_186 br_0_186 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c186
*+ bl_0_186 br_0_186 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c186
*+ bl_0_186 br_0_186 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c186
+ bl_0_186 br_0_186 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c187
+ bl_0_187 br_0_187 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c187
*+ bl_0_187 br_0_187 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c187
*+ bl_0_187 br_0_187 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c187
*+ bl_0_187 br_0_187 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c187
*+ bl_0_187 br_0_187 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c187
*+ bl_0_187 br_0_187 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c187
*+ bl_0_187 br_0_187 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c187
*+ bl_0_187 br_0_187 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c187
*+ bl_0_187 br_0_187 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c187
*+ bl_0_187 br_0_187 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c187
*+ bl_0_187 br_0_187 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c187
*+ bl_0_187 br_0_187 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c187
*+ bl_0_187 br_0_187 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c187
*+ bl_0_187 br_0_187 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c187
*+ bl_0_187 br_0_187 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c187
*+ bl_0_187 br_0_187 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c187
*+ bl_0_187 br_0_187 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c187
*+ bl_0_187 br_0_187 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c187
*+ bl_0_187 br_0_187 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c187
*+ bl_0_187 br_0_187 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c187
*+ bl_0_187 br_0_187 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c187
*+ bl_0_187 br_0_187 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c187
*+ bl_0_187 br_0_187 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c187
*+ bl_0_187 br_0_187 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c187
*+ bl_0_187 br_0_187 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c187
*+ bl_0_187 br_0_187 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c187
*+ bl_0_187 br_0_187 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c187
*+ bl_0_187 br_0_187 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c187
*+ bl_0_187 br_0_187 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c187
*+ bl_0_187 br_0_187 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c187
*+ bl_0_187 br_0_187 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c187
*+ bl_0_187 br_0_187 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c187
*+ bl_0_187 br_0_187 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c187
*+ bl_0_187 br_0_187 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c187
*+ bl_0_187 br_0_187 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c187
*+ bl_0_187 br_0_187 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c187
*+ bl_0_187 br_0_187 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c187
*+ bl_0_187 br_0_187 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c187
*+ bl_0_187 br_0_187 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c187
*+ bl_0_187 br_0_187 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c187
*+ bl_0_187 br_0_187 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c187
*+ bl_0_187 br_0_187 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c187
*+ bl_0_187 br_0_187 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c187
*+ bl_0_187 br_0_187 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c187
*+ bl_0_187 br_0_187 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c187
*+ bl_0_187 br_0_187 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c187
*+ bl_0_187 br_0_187 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c187
*+ bl_0_187 br_0_187 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c187
*+ bl_0_187 br_0_187 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c187
*+ bl_0_187 br_0_187 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c187
*+ bl_0_187 br_0_187 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c187
*+ bl_0_187 br_0_187 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c187
*+ bl_0_187 br_0_187 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c187
*+ bl_0_187 br_0_187 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c187
*+ bl_0_187 br_0_187 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c187
*+ bl_0_187 br_0_187 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c187
*+ bl_0_187 br_0_187 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c187
*+ bl_0_187 br_0_187 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c187
*+ bl_0_187 br_0_187 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c187
*+ bl_0_187 br_0_187 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c187
*+ bl_0_187 br_0_187 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c187
*+ bl_0_187 br_0_187 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c187
*+ bl_0_187 br_0_187 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c187
*+ bl_0_187 br_0_187 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c187
*+ bl_0_187 br_0_187 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c187
*+ bl_0_187 br_0_187 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c187
*+ bl_0_187 br_0_187 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c187
*+ bl_0_187 br_0_187 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c187
*+ bl_0_187 br_0_187 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c187
*+ bl_0_187 br_0_187 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c187
*+ bl_0_187 br_0_187 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c187
*+ bl_0_187 br_0_187 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c187
*+ bl_0_187 br_0_187 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c187
*+ bl_0_187 br_0_187 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c187
*+ bl_0_187 br_0_187 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c187
*+ bl_0_187 br_0_187 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c187
*+ bl_0_187 br_0_187 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c187
*+ bl_0_187 br_0_187 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c187
*+ bl_0_187 br_0_187 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c187
*+ bl_0_187 br_0_187 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c187
*+ bl_0_187 br_0_187 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c187
*+ bl_0_187 br_0_187 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c187
*+ bl_0_187 br_0_187 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c187
*+ bl_0_187 br_0_187 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c187
*+ bl_0_187 br_0_187 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c187
*+ bl_0_187 br_0_187 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c187
*+ bl_0_187 br_0_187 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c187
*+ bl_0_187 br_0_187 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c187
*+ bl_0_187 br_0_187 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c187
*+ bl_0_187 br_0_187 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c187
*+ bl_0_187 br_0_187 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c187
*+ bl_0_187 br_0_187 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c187
*+ bl_0_187 br_0_187 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c187
*+ bl_0_187 br_0_187 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c187
*+ bl_0_187 br_0_187 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c187
*+ bl_0_187 br_0_187 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c187
*+ bl_0_187 br_0_187 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c187
*+ bl_0_187 br_0_187 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c187
*+ bl_0_187 br_0_187 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c187
*+ bl_0_187 br_0_187 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c187
*+ bl_0_187 br_0_187 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c187
*+ bl_0_187 br_0_187 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c187
*+ bl_0_187 br_0_187 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c187
*+ bl_0_187 br_0_187 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c187
*+ bl_0_187 br_0_187 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c187
*+ bl_0_187 br_0_187 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c187
*+ bl_0_187 br_0_187 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c187
*+ bl_0_187 br_0_187 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c187
*+ bl_0_187 br_0_187 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c187
*+ bl_0_187 br_0_187 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c187
*+ bl_0_187 br_0_187 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c187
*+ bl_0_187 br_0_187 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c187
*+ bl_0_187 br_0_187 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c187
*+ bl_0_187 br_0_187 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c187
*+ bl_0_187 br_0_187 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c187
*+ bl_0_187 br_0_187 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c187
*+ bl_0_187 br_0_187 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c187
*+ bl_0_187 br_0_187 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c187
*+ bl_0_187 br_0_187 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c187
*+ bl_0_187 br_0_187 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c187
*+ bl_0_187 br_0_187 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c187
*+ bl_0_187 br_0_187 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c187
*+ bl_0_187 br_0_187 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c187
*+ bl_0_187 br_0_187 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c187
*+ bl_0_187 br_0_187 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c187
*+ bl_0_187 br_0_187 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c187
*+ bl_0_187 br_0_187 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c187
+ bl_0_187 br_0_187 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c188
+ bl_0_188 br_0_188 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c188
*+ bl_0_188 br_0_188 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c188
*+ bl_0_188 br_0_188 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c188
*+ bl_0_188 br_0_188 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c188
*+ bl_0_188 br_0_188 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c188
*+ bl_0_188 br_0_188 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c188
*+ bl_0_188 br_0_188 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c188
*+ bl_0_188 br_0_188 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c188
*+ bl_0_188 br_0_188 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c188
*+ bl_0_188 br_0_188 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c188
*+ bl_0_188 br_0_188 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c188
*+ bl_0_188 br_0_188 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c188
*+ bl_0_188 br_0_188 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c188
*+ bl_0_188 br_0_188 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c188
*+ bl_0_188 br_0_188 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c188
*+ bl_0_188 br_0_188 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c188
*+ bl_0_188 br_0_188 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c188
*+ bl_0_188 br_0_188 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c188
*+ bl_0_188 br_0_188 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c188
*+ bl_0_188 br_0_188 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c188
*+ bl_0_188 br_0_188 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c188
*+ bl_0_188 br_0_188 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c188
*+ bl_0_188 br_0_188 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c188
*+ bl_0_188 br_0_188 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c188
*+ bl_0_188 br_0_188 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c188
*+ bl_0_188 br_0_188 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c188
*+ bl_0_188 br_0_188 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c188
*+ bl_0_188 br_0_188 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c188
*+ bl_0_188 br_0_188 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c188
*+ bl_0_188 br_0_188 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c188
*+ bl_0_188 br_0_188 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c188
*+ bl_0_188 br_0_188 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c188
*+ bl_0_188 br_0_188 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c188
*+ bl_0_188 br_0_188 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c188
*+ bl_0_188 br_0_188 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c188
*+ bl_0_188 br_0_188 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c188
*+ bl_0_188 br_0_188 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c188
*+ bl_0_188 br_0_188 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c188
*+ bl_0_188 br_0_188 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c188
*+ bl_0_188 br_0_188 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c188
*+ bl_0_188 br_0_188 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c188
*+ bl_0_188 br_0_188 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c188
*+ bl_0_188 br_0_188 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c188
*+ bl_0_188 br_0_188 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c188
*+ bl_0_188 br_0_188 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c188
*+ bl_0_188 br_0_188 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c188
*+ bl_0_188 br_0_188 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c188
*+ bl_0_188 br_0_188 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c188
*+ bl_0_188 br_0_188 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c188
*+ bl_0_188 br_0_188 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c188
*+ bl_0_188 br_0_188 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c188
*+ bl_0_188 br_0_188 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c188
*+ bl_0_188 br_0_188 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c188
*+ bl_0_188 br_0_188 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c188
*+ bl_0_188 br_0_188 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c188
*+ bl_0_188 br_0_188 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c188
*+ bl_0_188 br_0_188 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c188
*+ bl_0_188 br_0_188 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c188
*+ bl_0_188 br_0_188 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c188
*+ bl_0_188 br_0_188 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c188
*+ bl_0_188 br_0_188 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c188
*+ bl_0_188 br_0_188 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c188
*+ bl_0_188 br_0_188 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c188
*+ bl_0_188 br_0_188 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c188
*+ bl_0_188 br_0_188 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c188
*+ bl_0_188 br_0_188 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c188
*+ bl_0_188 br_0_188 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c188
*+ bl_0_188 br_0_188 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c188
*+ bl_0_188 br_0_188 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c188
*+ bl_0_188 br_0_188 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c188
*+ bl_0_188 br_0_188 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c188
*+ bl_0_188 br_0_188 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c188
*+ bl_0_188 br_0_188 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c188
*+ bl_0_188 br_0_188 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c188
*+ bl_0_188 br_0_188 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c188
*+ bl_0_188 br_0_188 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c188
*+ bl_0_188 br_0_188 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c188
*+ bl_0_188 br_0_188 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c188
*+ bl_0_188 br_0_188 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c188
*+ bl_0_188 br_0_188 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c188
*+ bl_0_188 br_0_188 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c188
*+ bl_0_188 br_0_188 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c188
*+ bl_0_188 br_0_188 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c188
*+ bl_0_188 br_0_188 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c188
*+ bl_0_188 br_0_188 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c188
*+ bl_0_188 br_0_188 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c188
*+ bl_0_188 br_0_188 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c188
*+ bl_0_188 br_0_188 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c188
*+ bl_0_188 br_0_188 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c188
*+ bl_0_188 br_0_188 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c188
*+ bl_0_188 br_0_188 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c188
*+ bl_0_188 br_0_188 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c188
*+ bl_0_188 br_0_188 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c188
*+ bl_0_188 br_0_188 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c188
*+ bl_0_188 br_0_188 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c188
*+ bl_0_188 br_0_188 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c188
*+ bl_0_188 br_0_188 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c188
*+ bl_0_188 br_0_188 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c188
*+ bl_0_188 br_0_188 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c188
*+ bl_0_188 br_0_188 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c188
*+ bl_0_188 br_0_188 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c188
*+ bl_0_188 br_0_188 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c188
*+ bl_0_188 br_0_188 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c188
*+ bl_0_188 br_0_188 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c188
*+ bl_0_188 br_0_188 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c188
*+ bl_0_188 br_0_188 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c188
*+ bl_0_188 br_0_188 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c188
*+ bl_0_188 br_0_188 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c188
*+ bl_0_188 br_0_188 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c188
*+ bl_0_188 br_0_188 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c188
*+ bl_0_188 br_0_188 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c188
*+ bl_0_188 br_0_188 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c188
*+ bl_0_188 br_0_188 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c188
*+ bl_0_188 br_0_188 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c188
*+ bl_0_188 br_0_188 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c188
*+ bl_0_188 br_0_188 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c188
*+ bl_0_188 br_0_188 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c188
*+ bl_0_188 br_0_188 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c188
*+ bl_0_188 br_0_188 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c188
*+ bl_0_188 br_0_188 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c188
*+ bl_0_188 br_0_188 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c188
*+ bl_0_188 br_0_188 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c188
*+ bl_0_188 br_0_188 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c188
*+ bl_0_188 br_0_188 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c188
*+ bl_0_188 br_0_188 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c188
*+ bl_0_188 br_0_188 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c188
*+ bl_0_188 br_0_188 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c188
+ bl_0_188 br_0_188 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c189
+ bl_0_189 br_0_189 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c189
*+ bl_0_189 br_0_189 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c189
*+ bl_0_189 br_0_189 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c189
*+ bl_0_189 br_0_189 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c189
*+ bl_0_189 br_0_189 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c189
*+ bl_0_189 br_0_189 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c189
*+ bl_0_189 br_0_189 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c189
*+ bl_0_189 br_0_189 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c189
*+ bl_0_189 br_0_189 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c189
*+ bl_0_189 br_0_189 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c189
*+ bl_0_189 br_0_189 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c189
*+ bl_0_189 br_0_189 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c189
*+ bl_0_189 br_0_189 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c189
*+ bl_0_189 br_0_189 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c189
*+ bl_0_189 br_0_189 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c189
*+ bl_0_189 br_0_189 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c189
*+ bl_0_189 br_0_189 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c189
*+ bl_0_189 br_0_189 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c189
*+ bl_0_189 br_0_189 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c189
*+ bl_0_189 br_0_189 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c189
*+ bl_0_189 br_0_189 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c189
*+ bl_0_189 br_0_189 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c189
*+ bl_0_189 br_0_189 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c189
*+ bl_0_189 br_0_189 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c189
*+ bl_0_189 br_0_189 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c189
*+ bl_0_189 br_0_189 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c189
*+ bl_0_189 br_0_189 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c189
*+ bl_0_189 br_0_189 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c189
*+ bl_0_189 br_0_189 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c189
*+ bl_0_189 br_0_189 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c189
*+ bl_0_189 br_0_189 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c189
*+ bl_0_189 br_0_189 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c189
*+ bl_0_189 br_0_189 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c189
*+ bl_0_189 br_0_189 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c189
*+ bl_0_189 br_0_189 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c189
*+ bl_0_189 br_0_189 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c189
*+ bl_0_189 br_0_189 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c189
*+ bl_0_189 br_0_189 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c189
*+ bl_0_189 br_0_189 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c189
*+ bl_0_189 br_0_189 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c189
*+ bl_0_189 br_0_189 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c189
*+ bl_0_189 br_0_189 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c189
*+ bl_0_189 br_0_189 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c189
*+ bl_0_189 br_0_189 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c189
*+ bl_0_189 br_0_189 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c189
*+ bl_0_189 br_0_189 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c189
*+ bl_0_189 br_0_189 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c189
*+ bl_0_189 br_0_189 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c189
*+ bl_0_189 br_0_189 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c189
*+ bl_0_189 br_0_189 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c189
*+ bl_0_189 br_0_189 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c189
*+ bl_0_189 br_0_189 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c189
*+ bl_0_189 br_0_189 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c189
*+ bl_0_189 br_0_189 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c189
*+ bl_0_189 br_0_189 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c189
*+ bl_0_189 br_0_189 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c189
*+ bl_0_189 br_0_189 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c189
*+ bl_0_189 br_0_189 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c189
*+ bl_0_189 br_0_189 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c189
*+ bl_0_189 br_0_189 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c189
*+ bl_0_189 br_0_189 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c189
*+ bl_0_189 br_0_189 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c189
*+ bl_0_189 br_0_189 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c189
*+ bl_0_189 br_0_189 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c189
*+ bl_0_189 br_0_189 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c189
*+ bl_0_189 br_0_189 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c189
*+ bl_0_189 br_0_189 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c189
*+ bl_0_189 br_0_189 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c189
*+ bl_0_189 br_0_189 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c189
*+ bl_0_189 br_0_189 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c189
*+ bl_0_189 br_0_189 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c189
*+ bl_0_189 br_0_189 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c189
*+ bl_0_189 br_0_189 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c189
*+ bl_0_189 br_0_189 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c189
*+ bl_0_189 br_0_189 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c189
*+ bl_0_189 br_0_189 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c189
*+ bl_0_189 br_0_189 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c189
*+ bl_0_189 br_0_189 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c189
*+ bl_0_189 br_0_189 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c189
*+ bl_0_189 br_0_189 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c189
*+ bl_0_189 br_0_189 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c189
*+ bl_0_189 br_0_189 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c189
*+ bl_0_189 br_0_189 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c189
*+ bl_0_189 br_0_189 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c189
*+ bl_0_189 br_0_189 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c189
*+ bl_0_189 br_0_189 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c189
*+ bl_0_189 br_0_189 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c189
*+ bl_0_189 br_0_189 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c189
*+ bl_0_189 br_0_189 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c189
*+ bl_0_189 br_0_189 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c189
*+ bl_0_189 br_0_189 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c189
*+ bl_0_189 br_0_189 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c189
*+ bl_0_189 br_0_189 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c189
*+ bl_0_189 br_0_189 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c189
*+ bl_0_189 br_0_189 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c189
*+ bl_0_189 br_0_189 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c189
*+ bl_0_189 br_0_189 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c189
*+ bl_0_189 br_0_189 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c189
*+ bl_0_189 br_0_189 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c189
*+ bl_0_189 br_0_189 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c189
*+ bl_0_189 br_0_189 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c189
*+ bl_0_189 br_0_189 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c189
*+ bl_0_189 br_0_189 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c189
*+ bl_0_189 br_0_189 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c189
*+ bl_0_189 br_0_189 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c189
*+ bl_0_189 br_0_189 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c189
*+ bl_0_189 br_0_189 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c189
*+ bl_0_189 br_0_189 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c189
*+ bl_0_189 br_0_189 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c189
*+ bl_0_189 br_0_189 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c189
*+ bl_0_189 br_0_189 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c189
*+ bl_0_189 br_0_189 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c189
*+ bl_0_189 br_0_189 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c189
*+ bl_0_189 br_0_189 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c189
*+ bl_0_189 br_0_189 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c189
*+ bl_0_189 br_0_189 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c189
*+ bl_0_189 br_0_189 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c189
*+ bl_0_189 br_0_189 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c189
*+ bl_0_189 br_0_189 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c189
*+ bl_0_189 br_0_189 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c189
*+ bl_0_189 br_0_189 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c189
*+ bl_0_189 br_0_189 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c189
*+ bl_0_189 br_0_189 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c189
*+ bl_0_189 br_0_189 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c189
*+ bl_0_189 br_0_189 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c189
*+ bl_0_189 br_0_189 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c189
*+ bl_0_189 br_0_189 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c189
+ bl_0_189 br_0_189 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c190
+ bl_0_190 br_0_190 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c190
*+ bl_0_190 br_0_190 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c190
*+ bl_0_190 br_0_190 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c190
*+ bl_0_190 br_0_190 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c190
*+ bl_0_190 br_0_190 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c190
*+ bl_0_190 br_0_190 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c190
*+ bl_0_190 br_0_190 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c190
*+ bl_0_190 br_0_190 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c190
*+ bl_0_190 br_0_190 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c190
*+ bl_0_190 br_0_190 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c190
*+ bl_0_190 br_0_190 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c190
*+ bl_0_190 br_0_190 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c190
*+ bl_0_190 br_0_190 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c190
*+ bl_0_190 br_0_190 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c190
*+ bl_0_190 br_0_190 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c190
*+ bl_0_190 br_0_190 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c190
*+ bl_0_190 br_0_190 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c190
*+ bl_0_190 br_0_190 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c190
*+ bl_0_190 br_0_190 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c190
*+ bl_0_190 br_0_190 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c190
*+ bl_0_190 br_0_190 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c190
*+ bl_0_190 br_0_190 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c190
*+ bl_0_190 br_0_190 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c190
*+ bl_0_190 br_0_190 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c190
*+ bl_0_190 br_0_190 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c190
*+ bl_0_190 br_0_190 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c190
*+ bl_0_190 br_0_190 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c190
*+ bl_0_190 br_0_190 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c190
*+ bl_0_190 br_0_190 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c190
*+ bl_0_190 br_0_190 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c190
*+ bl_0_190 br_0_190 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c190
*+ bl_0_190 br_0_190 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c190
*+ bl_0_190 br_0_190 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c190
*+ bl_0_190 br_0_190 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c190
*+ bl_0_190 br_0_190 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c190
*+ bl_0_190 br_0_190 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c190
*+ bl_0_190 br_0_190 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c190
*+ bl_0_190 br_0_190 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c190
*+ bl_0_190 br_0_190 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c190
*+ bl_0_190 br_0_190 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c190
*+ bl_0_190 br_0_190 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c190
*+ bl_0_190 br_0_190 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c190
*+ bl_0_190 br_0_190 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c190
*+ bl_0_190 br_0_190 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c190
*+ bl_0_190 br_0_190 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c190
*+ bl_0_190 br_0_190 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c190
*+ bl_0_190 br_0_190 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c190
*+ bl_0_190 br_0_190 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c190
*+ bl_0_190 br_0_190 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c190
*+ bl_0_190 br_0_190 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c190
*+ bl_0_190 br_0_190 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c190
*+ bl_0_190 br_0_190 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c190
*+ bl_0_190 br_0_190 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c190
*+ bl_0_190 br_0_190 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c190
*+ bl_0_190 br_0_190 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c190
*+ bl_0_190 br_0_190 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c190
*+ bl_0_190 br_0_190 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c190
*+ bl_0_190 br_0_190 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c190
*+ bl_0_190 br_0_190 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c190
*+ bl_0_190 br_0_190 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c190
*+ bl_0_190 br_0_190 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c190
*+ bl_0_190 br_0_190 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c190
*+ bl_0_190 br_0_190 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c190
*+ bl_0_190 br_0_190 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c190
*+ bl_0_190 br_0_190 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c190
*+ bl_0_190 br_0_190 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c190
*+ bl_0_190 br_0_190 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c190
*+ bl_0_190 br_0_190 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c190
*+ bl_0_190 br_0_190 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c190
*+ bl_0_190 br_0_190 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c190
*+ bl_0_190 br_0_190 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c190
*+ bl_0_190 br_0_190 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c190
*+ bl_0_190 br_0_190 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c190
*+ bl_0_190 br_0_190 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c190
*+ bl_0_190 br_0_190 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c190
*+ bl_0_190 br_0_190 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c190
*+ bl_0_190 br_0_190 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c190
*+ bl_0_190 br_0_190 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c190
*+ bl_0_190 br_0_190 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c190
*+ bl_0_190 br_0_190 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c190
*+ bl_0_190 br_0_190 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c190
*+ bl_0_190 br_0_190 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c190
*+ bl_0_190 br_0_190 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c190
*+ bl_0_190 br_0_190 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c190
*+ bl_0_190 br_0_190 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c190
*+ bl_0_190 br_0_190 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c190
*+ bl_0_190 br_0_190 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c190
*+ bl_0_190 br_0_190 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c190
*+ bl_0_190 br_0_190 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c190
*+ bl_0_190 br_0_190 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c190
*+ bl_0_190 br_0_190 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c190
*+ bl_0_190 br_0_190 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c190
*+ bl_0_190 br_0_190 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c190
*+ bl_0_190 br_0_190 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c190
*+ bl_0_190 br_0_190 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c190
*+ bl_0_190 br_0_190 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c190
*+ bl_0_190 br_0_190 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c190
*+ bl_0_190 br_0_190 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c190
*+ bl_0_190 br_0_190 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c190
*+ bl_0_190 br_0_190 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c190
*+ bl_0_190 br_0_190 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c190
*+ bl_0_190 br_0_190 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c190
*+ bl_0_190 br_0_190 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c190
*+ bl_0_190 br_0_190 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c190
*+ bl_0_190 br_0_190 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c190
*+ bl_0_190 br_0_190 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c190
*+ bl_0_190 br_0_190 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c190
*+ bl_0_190 br_0_190 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c190
*+ bl_0_190 br_0_190 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c190
*+ bl_0_190 br_0_190 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c190
*+ bl_0_190 br_0_190 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c190
*+ bl_0_190 br_0_190 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c190
*+ bl_0_190 br_0_190 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c190
*+ bl_0_190 br_0_190 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c190
*+ bl_0_190 br_0_190 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c190
*+ bl_0_190 br_0_190 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c190
*+ bl_0_190 br_0_190 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c190
*+ bl_0_190 br_0_190 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c190
*+ bl_0_190 br_0_190 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c190
*+ bl_0_190 br_0_190 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c190
*+ bl_0_190 br_0_190 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c190
*+ bl_0_190 br_0_190 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c190
*+ bl_0_190 br_0_190 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c190
*+ bl_0_190 br_0_190 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c190
*+ bl_0_190 br_0_190 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c190
*+ bl_0_190 br_0_190 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c190
*+ bl_0_190 br_0_190 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c190
+ bl_0_190 br_0_190 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c191
+ bl_0_191 br_0_191 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c191
*+ bl_0_191 br_0_191 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c191
*+ bl_0_191 br_0_191 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c191
*+ bl_0_191 br_0_191 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c191
*+ bl_0_191 br_0_191 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c191
*+ bl_0_191 br_0_191 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c191
*+ bl_0_191 br_0_191 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c191
*+ bl_0_191 br_0_191 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c191
*+ bl_0_191 br_0_191 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c191
*+ bl_0_191 br_0_191 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c191
*+ bl_0_191 br_0_191 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c191
*+ bl_0_191 br_0_191 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c191
*+ bl_0_191 br_0_191 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c191
*+ bl_0_191 br_0_191 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c191
*+ bl_0_191 br_0_191 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c191
*+ bl_0_191 br_0_191 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c191
*+ bl_0_191 br_0_191 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c191
*+ bl_0_191 br_0_191 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c191
*+ bl_0_191 br_0_191 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c191
*+ bl_0_191 br_0_191 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c191
*+ bl_0_191 br_0_191 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c191
*+ bl_0_191 br_0_191 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c191
*+ bl_0_191 br_0_191 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c191
*+ bl_0_191 br_0_191 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c191
*+ bl_0_191 br_0_191 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c191
*+ bl_0_191 br_0_191 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c191
*+ bl_0_191 br_0_191 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c191
*+ bl_0_191 br_0_191 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c191
*+ bl_0_191 br_0_191 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c191
*+ bl_0_191 br_0_191 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c191
*+ bl_0_191 br_0_191 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c191
*+ bl_0_191 br_0_191 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c191
*+ bl_0_191 br_0_191 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c191
*+ bl_0_191 br_0_191 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c191
*+ bl_0_191 br_0_191 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c191
*+ bl_0_191 br_0_191 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c191
*+ bl_0_191 br_0_191 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c191
*+ bl_0_191 br_0_191 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c191
*+ bl_0_191 br_0_191 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c191
*+ bl_0_191 br_0_191 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c191
*+ bl_0_191 br_0_191 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c191
*+ bl_0_191 br_0_191 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c191
*+ bl_0_191 br_0_191 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c191
*+ bl_0_191 br_0_191 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c191
*+ bl_0_191 br_0_191 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c191
*+ bl_0_191 br_0_191 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c191
*+ bl_0_191 br_0_191 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c191
*+ bl_0_191 br_0_191 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c191
*+ bl_0_191 br_0_191 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c191
*+ bl_0_191 br_0_191 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c191
*+ bl_0_191 br_0_191 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c191
*+ bl_0_191 br_0_191 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c191
*+ bl_0_191 br_0_191 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c191
*+ bl_0_191 br_0_191 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c191
*+ bl_0_191 br_0_191 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c191
*+ bl_0_191 br_0_191 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c191
*+ bl_0_191 br_0_191 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c191
*+ bl_0_191 br_0_191 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c191
*+ bl_0_191 br_0_191 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c191
*+ bl_0_191 br_0_191 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c191
*+ bl_0_191 br_0_191 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c191
*+ bl_0_191 br_0_191 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c191
*+ bl_0_191 br_0_191 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c191
*+ bl_0_191 br_0_191 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c191
*+ bl_0_191 br_0_191 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c191
*+ bl_0_191 br_0_191 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c191
*+ bl_0_191 br_0_191 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c191
*+ bl_0_191 br_0_191 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c191
*+ bl_0_191 br_0_191 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c191
*+ bl_0_191 br_0_191 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c191
*+ bl_0_191 br_0_191 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c191
*+ bl_0_191 br_0_191 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c191
*+ bl_0_191 br_0_191 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c191
*+ bl_0_191 br_0_191 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c191
*+ bl_0_191 br_0_191 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c191
*+ bl_0_191 br_0_191 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c191
*+ bl_0_191 br_0_191 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c191
*+ bl_0_191 br_0_191 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c191
*+ bl_0_191 br_0_191 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c191
*+ bl_0_191 br_0_191 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c191
*+ bl_0_191 br_0_191 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c191
*+ bl_0_191 br_0_191 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c191
*+ bl_0_191 br_0_191 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c191
*+ bl_0_191 br_0_191 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c191
*+ bl_0_191 br_0_191 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c191
*+ bl_0_191 br_0_191 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c191
*+ bl_0_191 br_0_191 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c191
*+ bl_0_191 br_0_191 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c191
*+ bl_0_191 br_0_191 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c191
*+ bl_0_191 br_0_191 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c191
*+ bl_0_191 br_0_191 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c191
*+ bl_0_191 br_0_191 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c191
*+ bl_0_191 br_0_191 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c191
*+ bl_0_191 br_0_191 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c191
*+ bl_0_191 br_0_191 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c191
*+ bl_0_191 br_0_191 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c191
*+ bl_0_191 br_0_191 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c191
*+ bl_0_191 br_0_191 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c191
*+ bl_0_191 br_0_191 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c191
*+ bl_0_191 br_0_191 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c191
*+ bl_0_191 br_0_191 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c191
*+ bl_0_191 br_0_191 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c191
*+ bl_0_191 br_0_191 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c191
*+ bl_0_191 br_0_191 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c191
*+ bl_0_191 br_0_191 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c191
*+ bl_0_191 br_0_191 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c191
*+ bl_0_191 br_0_191 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c191
*+ bl_0_191 br_0_191 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c191
*+ bl_0_191 br_0_191 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c191
*+ bl_0_191 br_0_191 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c191
*+ bl_0_191 br_0_191 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c191
*+ bl_0_191 br_0_191 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c191
*+ bl_0_191 br_0_191 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c191
*+ bl_0_191 br_0_191 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c191
*+ bl_0_191 br_0_191 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c191
*+ bl_0_191 br_0_191 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c191
*+ bl_0_191 br_0_191 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c191
*+ bl_0_191 br_0_191 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c191
*+ bl_0_191 br_0_191 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c191
*+ bl_0_191 br_0_191 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c191
*+ bl_0_191 br_0_191 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c191
*+ bl_0_191 br_0_191 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c191
*+ bl_0_191 br_0_191 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c191
*+ bl_0_191 br_0_191 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c191
*+ bl_0_191 br_0_191 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c191
*+ bl_0_191 br_0_191 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c191
*+ bl_0_191 br_0_191 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c191
+ bl_0_191 br_0_191 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c192
+ bl_0_192 br_0_192 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c192
*+ bl_0_192 br_0_192 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c192
*+ bl_0_192 br_0_192 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c192
*+ bl_0_192 br_0_192 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c192
*+ bl_0_192 br_0_192 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c192
*+ bl_0_192 br_0_192 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c192
*+ bl_0_192 br_0_192 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c192
*+ bl_0_192 br_0_192 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c192
*+ bl_0_192 br_0_192 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c192
*+ bl_0_192 br_0_192 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c192
*+ bl_0_192 br_0_192 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c192
*+ bl_0_192 br_0_192 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c192
*+ bl_0_192 br_0_192 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c192
*+ bl_0_192 br_0_192 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c192
*+ bl_0_192 br_0_192 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c192
*+ bl_0_192 br_0_192 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c192
*+ bl_0_192 br_0_192 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c192
*+ bl_0_192 br_0_192 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c192
*+ bl_0_192 br_0_192 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c192
*+ bl_0_192 br_0_192 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c192
*+ bl_0_192 br_0_192 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c192
*+ bl_0_192 br_0_192 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c192
*+ bl_0_192 br_0_192 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c192
*+ bl_0_192 br_0_192 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c192
*+ bl_0_192 br_0_192 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c192
*+ bl_0_192 br_0_192 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c192
*+ bl_0_192 br_0_192 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c192
*+ bl_0_192 br_0_192 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c192
*+ bl_0_192 br_0_192 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c192
*+ bl_0_192 br_0_192 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c192
*+ bl_0_192 br_0_192 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c192
*+ bl_0_192 br_0_192 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c192
*+ bl_0_192 br_0_192 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c192
*+ bl_0_192 br_0_192 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c192
*+ bl_0_192 br_0_192 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c192
*+ bl_0_192 br_0_192 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c192
*+ bl_0_192 br_0_192 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c192
*+ bl_0_192 br_0_192 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c192
*+ bl_0_192 br_0_192 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c192
*+ bl_0_192 br_0_192 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c192
*+ bl_0_192 br_0_192 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c192
*+ bl_0_192 br_0_192 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c192
*+ bl_0_192 br_0_192 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c192
*+ bl_0_192 br_0_192 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c192
*+ bl_0_192 br_0_192 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c192
*+ bl_0_192 br_0_192 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c192
*+ bl_0_192 br_0_192 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c192
*+ bl_0_192 br_0_192 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c192
*+ bl_0_192 br_0_192 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c192
*+ bl_0_192 br_0_192 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c192
*+ bl_0_192 br_0_192 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c192
*+ bl_0_192 br_0_192 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c192
*+ bl_0_192 br_0_192 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c192
*+ bl_0_192 br_0_192 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c192
*+ bl_0_192 br_0_192 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c192
*+ bl_0_192 br_0_192 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c192
*+ bl_0_192 br_0_192 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c192
*+ bl_0_192 br_0_192 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c192
*+ bl_0_192 br_0_192 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c192
*+ bl_0_192 br_0_192 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c192
*+ bl_0_192 br_0_192 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c192
*+ bl_0_192 br_0_192 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c192
*+ bl_0_192 br_0_192 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c192
*+ bl_0_192 br_0_192 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c192
*+ bl_0_192 br_0_192 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c192
*+ bl_0_192 br_0_192 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c192
*+ bl_0_192 br_0_192 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c192
*+ bl_0_192 br_0_192 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c192
*+ bl_0_192 br_0_192 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c192
*+ bl_0_192 br_0_192 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c192
*+ bl_0_192 br_0_192 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c192
*+ bl_0_192 br_0_192 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c192
*+ bl_0_192 br_0_192 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c192
*+ bl_0_192 br_0_192 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c192
*+ bl_0_192 br_0_192 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c192
*+ bl_0_192 br_0_192 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c192
*+ bl_0_192 br_0_192 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c192
*+ bl_0_192 br_0_192 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c192
*+ bl_0_192 br_0_192 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c192
*+ bl_0_192 br_0_192 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c192
*+ bl_0_192 br_0_192 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c192
*+ bl_0_192 br_0_192 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c192
*+ bl_0_192 br_0_192 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c192
*+ bl_0_192 br_0_192 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c192
*+ bl_0_192 br_0_192 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c192
*+ bl_0_192 br_0_192 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c192
*+ bl_0_192 br_0_192 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c192
*+ bl_0_192 br_0_192 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c192
*+ bl_0_192 br_0_192 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c192
*+ bl_0_192 br_0_192 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c192
*+ bl_0_192 br_0_192 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c192
*+ bl_0_192 br_0_192 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c192
*+ bl_0_192 br_0_192 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c192
*+ bl_0_192 br_0_192 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c192
*+ bl_0_192 br_0_192 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c192
*+ bl_0_192 br_0_192 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c192
*+ bl_0_192 br_0_192 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c192
*+ bl_0_192 br_0_192 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c192
*+ bl_0_192 br_0_192 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c192
*+ bl_0_192 br_0_192 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c192
*+ bl_0_192 br_0_192 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c192
*+ bl_0_192 br_0_192 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c192
*+ bl_0_192 br_0_192 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c192
*+ bl_0_192 br_0_192 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c192
*+ bl_0_192 br_0_192 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c192
*+ bl_0_192 br_0_192 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c192
*+ bl_0_192 br_0_192 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c192
*+ bl_0_192 br_0_192 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c192
*+ bl_0_192 br_0_192 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c192
*+ bl_0_192 br_0_192 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c192
*+ bl_0_192 br_0_192 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c192
*+ bl_0_192 br_0_192 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c192
*+ bl_0_192 br_0_192 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c192
*+ bl_0_192 br_0_192 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c192
*+ bl_0_192 br_0_192 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c192
*+ bl_0_192 br_0_192 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c192
*+ bl_0_192 br_0_192 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c192
*+ bl_0_192 br_0_192 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c192
*+ bl_0_192 br_0_192 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c192
*+ bl_0_192 br_0_192 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c192
*+ bl_0_192 br_0_192 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c192
*+ bl_0_192 br_0_192 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c192
*+ bl_0_192 br_0_192 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c192
*+ bl_0_192 br_0_192 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c192
*+ bl_0_192 br_0_192 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c192
*+ bl_0_192 br_0_192 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c192
*+ bl_0_192 br_0_192 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c192
+ bl_0_192 br_0_192 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c193
+ bl_0_193 br_0_193 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c193
*+ bl_0_193 br_0_193 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c193
*+ bl_0_193 br_0_193 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c193
*+ bl_0_193 br_0_193 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c193
*+ bl_0_193 br_0_193 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c193
*+ bl_0_193 br_0_193 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c193
*+ bl_0_193 br_0_193 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c193
*+ bl_0_193 br_0_193 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c193
*+ bl_0_193 br_0_193 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c193
*+ bl_0_193 br_0_193 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c193
*+ bl_0_193 br_0_193 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c193
*+ bl_0_193 br_0_193 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c193
*+ bl_0_193 br_0_193 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c193
*+ bl_0_193 br_0_193 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c193
*+ bl_0_193 br_0_193 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c193
*+ bl_0_193 br_0_193 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c193
*+ bl_0_193 br_0_193 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c193
*+ bl_0_193 br_0_193 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c193
*+ bl_0_193 br_0_193 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c193
*+ bl_0_193 br_0_193 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c193
*+ bl_0_193 br_0_193 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c193
*+ bl_0_193 br_0_193 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c193
*+ bl_0_193 br_0_193 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c193
*+ bl_0_193 br_0_193 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c193
*+ bl_0_193 br_0_193 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c193
*+ bl_0_193 br_0_193 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c193
*+ bl_0_193 br_0_193 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c193
*+ bl_0_193 br_0_193 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c193
*+ bl_0_193 br_0_193 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c193
*+ bl_0_193 br_0_193 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c193
*+ bl_0_193 br_0_193 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c193
*+ bl_0_193 br_0_193 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c193
*+ bl_0_193 br_0_193 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c193
*+ bl_0_193 br_0_193 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c193
*+ bl_0_193 br_0_193 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c193
*+ bl_0_193 br_0_193 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c193
*+ bl_0_193 br_0_193 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c193
*+ bl_0_193 br_0_193 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c193
*+ bl_0_193 br_0_193 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c193
*+ bl_0_193 br_0_193 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c193
*+ bl_0_193 br_0_193 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c193
*+ bl_0_193 br_0_193 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c193
*+ bl_0_193 br_0_193 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c193
*+ bl_0_193 br_0_193 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c193
*+ bl_0_193 br_0_193 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c193
*+ bl_0_193 br_0_193 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c193
*+ bl_0_193 br_0_193 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c193
*+ bl_0_193 br_0_193 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c193
*+ bl_0_193 br_0_193 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c193
*+ bl_0_193 br_0_193 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c193
*+ bl_0_193 br_0_193 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c193
*+ bl_0_193 br_0_193 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c193
*+ bl_0_193 br_0_193 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c193
*+ bl_0_193 br_0_193 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c193
*+ bl_0_193 br_0_193 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c193
*+ bl_0_193 br_0_193 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c193
*+ bl_0_193 br_0_193 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c193
*+ bl_0_193 br_0_193 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c193
*+ bl_0_193 br_0_193 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c193
*+ bl_0_193 br_0_193 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c193
*+ bl_0_193 br_0_193 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c193
*+ bl_0_193 br_0_193 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c193
*+ bl_0_193 br_0_193 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c193
*+ bl_0_193 br_0_193 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c193
*+ bl_0_193 br_0_193 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c193
*+ bl_0_193 br_0_193 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c193
*+ bl_0_193 br_0_193 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c193
*+ bl_0_193 br_0_193 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c193
*+ bl_0_193 br_0_193 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c193
*+ bl_0_193 br_0_193 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c193
*+ bl_0_193 br_0_193 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c193
*+ bl_0_193 br_0_193 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c193
*+ bl_0_193 br_0_193 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c193
*+ bl_0_193 br_0_193 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c193
*+ bl_0_193 br_0_193 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c193
*+ bl_0_193 br_0_193 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c193
*+ bl_0_193 br_0_193 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c193
*+ bl_0_193 br_0_193 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c193
*+ bl_0_193 br_0_193 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c193
*+ bl_0_193 br_0_193 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c193
*+ bl_0_193 br_0_193 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c193
*+ bl_0_193 br_0_193 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c193
*+ bl_0_193 br_0_193 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c193
*+ bl_0_193 br_0_193 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c193
*+ bl_0_193 br_0_193 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c193
*+ bl_0_193 br_0_193 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c193
*+ bl_0_193 br_0_193 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c193
*+ bl_0_193 br_0_193 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c193
*+ bl_0_193 br_0_193 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c193
*+ bl_0_193 br_0_193 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c193
*+ bl_0_193 br_0_193 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c193
*+ bl_0_193 br_0_193 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c193
*+ bl_0_193 br_0_193 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c193
*+ bl_0_193 br_0_193 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c193
*+ bl_0_193 br_0_193 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c193
*+ bl_0_193 br_0_193 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c193
*+ bl_0_193 br_0_193 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c193
*+ bl_0_193 br_0_193 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c193
*+ bl_0_193 br_0_193 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c193
*+ bl_0_193 br_0_193 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c193
*+ bl_0_193 br_0_193 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c193
*+ bl_0_193 br_0_193 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c193
*+ bl_0_193 br_0_193 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c193
*+ bl_0_193 br_0_193 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c193
*+ bl_0_193 br_0_193 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c193
*+ bl_0_193 br_0_193 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c193
*+ bl_0_193 br_0_193 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c193
*+ bl_0_193 br_0_193 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c193
*+ bl_0_193 br_0_193 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c193
*+ bl_0_193 br_0_193 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c193
*+ bl_0_193 br_0_193 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c193
*+ bl_0_193 br_0_193 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c193
*+ bl_0_193 br_0_193 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c193
*+ bl_0_193 br_0_193 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c193
*+ bl_0_193 br_0_193 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c193
*+ bl_0_193 br_0_193 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c193
*+ bl_0_193 br_0_193 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c193
*+ bl_0_193 br_0_193 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c193
*+ bl_0_193 br_0_193 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c193
*+ bl_0_193 br_0_193 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c193
*+ bl_0_193 br_0_193 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c193
*+ bl_0_193 br_0_193 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c193
*+ bl_0_193 br_0_193 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c193
*+ bl_0_193 br_0_193 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c193
*+ bl_0_193 br_0_193 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c193
*+ bl_0_193 br_0_193 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c193
*+ bl_0_193 br_0_193 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c193
+ bl_0_193 br_0_193 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c194
+ bl_0_194 br_0_194 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c194
*+ bl_0_194 br_0_194 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c194
*+ bl_0_194 br_0_194 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c194
*+ bl_0_194 br_0_194 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c194
*+ bl_0_194 br_0_194 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c194
*+ bl_0_194 br_0_194 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c194
*+ bl_0_194 br_0_194 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c194
*+ bl_0_194 br_0_194 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c194
*+ bl_0_194 br_0_194 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c194
*+ bl_0_194 br_0_194 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c194
*+ bl_0_194 br_0_194 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c194
*+ bl_0_194 br_0_194 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c194
*+ bl_0_194 br_0_194 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c194
*+ bl_0_194 br_0_194 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c194
*+ bl_0_194 br_0_194 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c194
*+ bl_0_194 br_0_194 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c194
*+ bl_0_194 br_0_194 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c194
*+ bl_0_194 br_0_194 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c194
*+ bl_0_194 br_0_194 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c194
*+ bl_0_194 br_0_194 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c194
*+ bl_0_194 br_0_194 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c194
*+ bl_0_194 br_0_194 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c194
*+ bl_0_194 br_0_194 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c194
*+ bl_0_194 br_0_194 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c194
*+ bl_0_194 br_0_194 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c194
*+ bl_0_194 br_0_194 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c194
*+ bl_0_194 br_0_194 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c194
*+ bl_0_194 br_0_194 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c194
*+ bl_0_194 br_0_194 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c194
*+ bl_0_194 br_0_194 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c194
*+ bl_0_194 br_0_194 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c194
*+ bl_0_194 br_0_194 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c194
*+ bl_0_194 br_0_194 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c194
*+ bl_0_194 br_0_194 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c194
*+ bl_0_194 br_0_194 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c194
*+ bl_0_194 br_0_194 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c194
*+ bl_0_194 br_0_194 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c194
*+ bl_0_194 br_0_194 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c194
*+ bl_0_194 br_0_194 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c194
*+ bl_0_194 br_0_194 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c194
*+ bl_0_194 br_0_194 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c194
*+ bl_0_194 br_0_194 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c194
*+ bl_0_194 br_0_194 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c194
*+ bl_0_194 br_0_194 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c194
*+ bl_0_194 br_0_194 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c194
*+ bl_0_194 br_0_194 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c194
*+ bl_0_194 br_0_194 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c194
*+ bl_0_194 br_0_194 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c194
*+ bl_0_194 br_0_194 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c194
*+ bl_0_194 br_0_194 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c194
*+ bl_0_194 br_0_194 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c194
*+ bl_0_194 br_0_194 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c194
*+ bl_0_194 br_0_194 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c194
*+ bl_0_194 br_0_194 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c194
*+ bl_0_194 br_0_194 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c194
*+ bl_0_194 br_0_194 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c194
*+ bl_0_194 br_0_194 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c194
*+ bl_0_194 br_0_194 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c194
*+ bl_0_194 br_0_194 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c194
*+ bl_0_194 br_0_194 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c194
*+ bl_0_194 br_0_194 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c194
*+ bl_0_194 br_0_194 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c194
*+ bl_0_194 br_0_194 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c194
*+ bl_0_194 br_0_194 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c194
*+ bl_0_194 br_0_194 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c194
*+ bl_0_194 br_0_194 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c194
*+ bl_0_194 br_0_194 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c194
*+ bl_0_194 br_0_194 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c194
*+ bl_0_194 br_0_194 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c194
*+ bl_0_194 br_0_194 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c194
*+ bl_0_194 br_0_194 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c194
*+ bl_0_194 br_0_194 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c194
*+ bl_0_194 br_0_194 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c194
*+ bl_0_194 br_0_194 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c194
*+ bl_0_194 br_0_194 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c194
*+ bl_0_194 br_0_194 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c194
*+ bl_0_194 br_0_194 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c194
*+ bl_0_194 br_0_194 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c194
*+ bl_0_194 br_0_194 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c194
*+ bl_0_194 br_0_194 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c194
*+ bl_0_194 br_0_194 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c194
*+ bl_0_194 br_0_194 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c194
*+ bl_0_194 br_0_194 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c194
*+ bl_0_194 br_0_194 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c194
*+ bl_0_194 br_0_194 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c194
*+ bl_0_194 br_0_194 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c194
*+ bl_0_194 br_0_194 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c194
*+ bl_0_194 br_0_194 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c194
*+ bl_0_194 br_0_194 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c194
*+ bl_0_194 br_0_194 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c194
*+ bl_0_194 br_0_194 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c194
*+ bl_0_194 br_0_194 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c194
*+ bl_0_194 br_0_194 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c194
*+ bl_0_194 br_0_194 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c194
*+ bl_0_194 br_0_194 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c194
*+ bl_0_194 br_0_194 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c194
*+ bl_0_194 br_0_194 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c194
*+ bl_0_194 br_0_194 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c194
*+ bl_0_194 br_0_194 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c194
*+ bl_0_194 br_0_194 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c194
*+ bl_0_194 br_0_194 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c194
*+ bl_0_194 br_0_194 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c194
*+ bl_0_194 br_0_194 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c194
*+ bl_0_194 br_0_194 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c194
*+ bl_0_194 br_0_194 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c194
*+ bl_0_194 br_0_194 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c194
*+ bl_0_194 br_0_194 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c194
*+ bl_0_194 br_0_194 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c194
*+ bl_0_194 br_0_194 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c194
*+ bl_0_194 br_0_194 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c194
*+ bl_0_194 br_0_194 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c194
*+ bl_0_194 br_0_194 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c194
*+ bl_0_194 br_0_194 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c194
*+ bl_0_194 br_0_194 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c194
*+ bl_0_194 br_0_194 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c194
*+ bl_0_194 br_0_194 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c194
*+ bl_0_194 br_0_194 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c194
*+ bl_0_194 br_0_194 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c194
*+ bl_0_194 br_0_194 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c194
*+ bl_0_194 br_0_194 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c194
*+ bl_0_194 br_0_194 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c194
*+ bl_0_194 br_0_194 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c194
*+ bl_0_194 br_0_194 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c194
*+ bl_0_194 br_0_194 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c194
*+ bl_0_194 br_0_194 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c194
*+ bl_0_194 br_0_194 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c194
*+ bl_0_194 br_0_194 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c194
+ bl_0_194 br_0_194 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c195
+ bl_0_195 br_0_195 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c195
*+ bl_0_195 br_0_195 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c195
*+ bl_0_195 br_0_195 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c195
*+ bl_0_195 br_0_195 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c195
*+ bl_0_195 br_0_195 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c195
*+ bl_0_195 br_0_195 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c195
*+ bl_0_195 br_0_195 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c195
*+ bl_0_195 br_0_195 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c195
*+ bl_0_195 br_0_195 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c195
*+ bl_0_195 br_0_195 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c195
*+ bl_0_195 br_0_195 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c195
*+ bl_0_195 br_0_195 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c195
*+ bl_0_195 br_0_195 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c195
*+ bl_0_195 br_0_195 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c195
*+ bl_0_195 br_0_195 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c195
*+ bl_0_195 br_0_195 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c195
*+ bl_0_195 br_0_195 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c195
*+ bl_0_195 br_0_195 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c195
*+ bl_0_195 br_0_195 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c195
*+ bl_0_195 br_0_195 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c195
*+ bl_0_195 br_0_195 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c195
*+ bl_0_195 br_0_195 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c195
*+ bl_0_195 br_0_195 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c195
*+ bl_0_195 br_0_195 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c195
*+ bl_0_195 br_0_195 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c195
*+ bl_0_195 br_0_195 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c195
*+ bl_0_195 br_0_195 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c195
*+ bl_0_195 br_0_195 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c195
*+ bl_0_195 br_0_195 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c195
*+ bl_0_195 br_0_195 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c195
*+ bl_0_195 br_0_195 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c195
*+ bl_0_195 br_0_195 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c195
*+ bl_0_195 br_0_195 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c195
*+ bl_0_195 br_0_195 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c195
*+ bl_0_195 br_0_195 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c195
*+ bl_0_195 br_0_195 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c195
*+ bl_0_195 br_0_195 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c195
*+ bl_0_195 br_0_195 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c195
*+ bl_0_195 br_0_195 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c195
*+ bl_0_195 br_0_195 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c195
*+ bl_0_195 br_0_195 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c195
*+ bl_0_195 br_0_195 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c195
*+ bl_0_195 br_0_195 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c195
*+ bl_0_195 br_0_195 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c195
*+ bl_0_195 br_0_195 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c195
*+ bl_0_195 br_0_195 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c195
*+ bl_0_195 br_0_195 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c195
*+ bl_0_195 br_0_195 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c195
*+ bl_0_195 br_0_195 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c195
*+ bl_0_195 br_0_195 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c195
*+ bl_0_195 br_0_195 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c195
*+ bl_0_195 br_0_195 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c195
*+ bl_0_195 br_0_195 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c195
*+ bl_0_195 br_0_195 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c195
*+ bl_0_195 br_0_195 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c195
*+ bl_0_195 br_0_195 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c195
*+ bl_0_195 br_0_195 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c195
*+ bl_0_195 br_0_195 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c195
*+ bl_0_195 br_0_195 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c195
*+ bl_0_195 br_0_195 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c195
*+ bl_0_195 br_0_195 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c195
*+ bl_0_195 br_0_195 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c195
*+ bl_0_195 br_0_195 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c195
*+ bl_0_195 br_0_195 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c195
*+ bl_0_195 br_0_195 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c195
*+ bl_0_195 br_0_195 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c195
*+ bl_0_195 br_0_195 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c195
*+ bl_0_195 br_0_195 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c195
*+ bl_0_195 br_0_195 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c195
*+ bl_0_195 br_0_195 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c195
*+ bl_0_195 br_0_195 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c195
*+ bl_0_195 br_0_195 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c195
*+ bl_0_195 br_0_195 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c195
*+ bl_0_195 br_0_195 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c195
*+ bl_0_195 br_0_195 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c195
*+ bl_0_195 br_0_195 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c195
*+ bl_0_195 br_0_195 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c195
*+ bl_0_195 br_0_195 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c195
*+ bl_0_195 br_0_195 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c195
*+ bl_0_195 br_0_195 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c195
*+ bl_0_195 br_0_195 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c195
*+ bl_0_195 br_0_195 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c195
*+ bl_0_195 br_0_195 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c195
*+ bl_0_195 br_0_195 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c195
*+ bl_0_195 br_0_195 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c195
*+ bl_0_195 br_0_195 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c195
*+ bl_0_195 br_0_195 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c195
*+ bl_0_195 br_0_195 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c195
*+ bl_0_195 br_0_195 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c195
*+ bl_0_195 br_0_195 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c195
*+ bl_0_195 br_0_195 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c195
*+ bl_0_195 br_0_195 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c195
*+ bl_0_195 br_0_195 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c195
*+ bl_0_195 br_0_195 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c195
*+ bl_0_195 br_0_195 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c195
*+ bl_0_195 br_0_195 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c195
*+ bl_0_195 br_0_195 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c195
*+ bl_0_195 br_0_195 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c195
*+ bl_0_195 br_0_195 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c195
*+ bl_0_195 br_0_195 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c195
*+ bl_0_195 br_0_195 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c195
*+ bl_0_195 br_0_195 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c195
*+ bl_0_195 br_0_195 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c195
*+ bl_0_195 br_0_195 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c195
*+ bl_0_195 br_0_195 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c195
*+ bl_0_195 br_0_195 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c195
*+ bl_0_195 br_0_195 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c195
*+ bl_0_195 br_0_195 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c195
*+ bl_0_195 br_0_195 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c195
*+ bl_0_195 br_0_195 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c195
*+ bl_0_195 br_0_195 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c195
*+ bl_0_195 br_0_195 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c195
*+ bl_0_195 br_0_195 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c195
*+ bl_0_195 br_0_195 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c195
*+ bl_0_195 br_0_195 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c195
*+ bl_0_195 br_0_195 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c195
*+ bl_0_195 br_0_195 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c195
*+ bl_0_195 br_0_195 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c195
*+ bl_0_195 br_0_195 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c195
*+ bl_0_195 br_0_195 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c195
*+ bl_0_195 br_0_195 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c195
*+ bl_0_195 br_0_195 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c195
*+ bl_0_195 br_0_195 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c195
*+ bl_0_195 br_0_195 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c195
*+ bl_0_195 br_0_195 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c195
*+ bl_0_195 br_0_195 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c195
*+ bl_0_195 br_0_195 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c195
+ bl_0_195 br_0_195 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c196
+ bl_0_196 br_0_196 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c196
*+ bl_0_196 br_0_196 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c196
*+ bl_0_196 br_0_196 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c196
*+ bl_0_196 br_0_196 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c196
*+ bl_0_196 br_0_196 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c196
*+ bl_0_196 br_0_196 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c196
*+ bl_0_196 br_0_196 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c196
*+ bl_0_196 br_0_196 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c196
*+ bl_0_196 br_0_196 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c196
*+ bl_0_196 br_0_196 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c196
*+ bl_0_196 br_0_196 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c196
*+ bl_0_196 br_0_196 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c196
*+ bl_0_196 br_0_196 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c196
*+ bl_0_196 br_0_196 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c196
*+ bl_0_196 br_0_196 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c196
*+ bl_0_196 br_0_196 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c196
*+ bl_0_196 br_0_196 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c196
*+ bl_0_196 br_0_196 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c196
*+ bl_0_196 br_0_196 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c196
*+ bl_0_196 br_0_196 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c196
*+ bl_0_196 br_0_196 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c196
*+ bl_0_196 br_0_196 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c196
*+ bl_0_196 br_0_196 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c196
*+ bl_0_196 br_0_196 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c196
*+ bl_0_196 br_0_196 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c196
*+ bl_0_196 br_0_196 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c196
*+ bl_0_196 br_0_196 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c196
*+ bl_0_196 br_0_196 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c196
*+ bl_0_196 br_0_196 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c196
*+ bl_0_196 br_0_196 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c196
*+ bl_0_196 br_0_196 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c196
*+ bl_0_196 br_0_196 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c196
*+ bl_0_196 br_0_196 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c196
*+ bl_0_196 br_0_196 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c196
*+ bl_0_196 br_0_196 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c196
*+ bl_0_196 br_0_196 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c196
*+ bl_0_196 br_0_196 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c196
*+ bl_0_196 br_0_196 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c196
*+ bl_0_196 br_0_196 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c196
*+ bl_0_196 br_0_196 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c196
*+ bl_0_196 br_0_196 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c196
*+ bl_0_196 br_0_196 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c196
*+ bl_0_196 br_0_196 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c196
*+ bl_0_196 br_0_196 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c196
*+ bl_0_196 br_0_196 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c196
*+ bl_0_196 br_0_196 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c196
*+ bl_0_196 br_0_196 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c196
*+ bl_0_196 br_0_196 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c196
*+ bl_0_196 br_0_196 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c196
*+ bl_0_196 br_0_196 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c196
*+ bl_0_196 br_0_196 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c196
*+ bl_0_196 br_0_196 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c196
*+ bl_0_196 br_0_196 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c196
*+ bl_0_196 br_0_196 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c196
*+ bl_0_196 br_0_196 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c196
*+ bl_0_196 br_0_196 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c196
*+ bl_0_196 br_0_196 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c196
*+ bl_0_196 br_0_196 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c196
*+ bl_0_196 br_0_196 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c196
*+ bl_0_196 br_0_196 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c196
*+ bl_0_196 br_0_196 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c196
*+ bl_0_196 br_0_196 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c196
*+ bl_0_196 br_0_196 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c196
*+ bl_0_196 br_0_196 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c196
*+ bl_0_196 br_0_196 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c196
*+ bl_0_196 br_0_196 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c196
*+ bl_0_196 br_0_196 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c196
*+ bl_0_196 br_0_196 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c196
*+ bl_0_196 br_0_196 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c196
*+ bl_0_196 br_0_196 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c196
*+ bl_0_196 br_0_196 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c196
*+ bl_0_196 br_0_196 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c196
*+ bl_0_196 br_0_196 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c196
*+ bl_0_196 br_0_196 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c196
*+ bl_0_196 br_0_196 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c196
*+ bl_0_196 br_0_196 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c196
*+ bl_0_196 br_0_196 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c196
*+ bl_0_196 br_0_196 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c196
*+ bl_0_196 br_0_196 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c196
*+ bl_0_196 br_0_196 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c196
*+ bl_0_196 br_0_196 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c196
*+ bl_0_196 br_0_196 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c196
*+ bl_0_196 br_0_196 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c196
*+ bl_0_196 br_0_196 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c196
*+ bl_0_196 br_0_196 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c196
*+ bl_0_196 br_0_196 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c196
*+ bl_0_196 br_0_196 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c196
*+ bl_0_196 br_0_196 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c196
*+ bl_0_196 br_0_196 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c196
*+ bl_0_196 br_0_196 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c196
*+ bl_0_196 br_0_196 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c196
*+ bl_0_196 br_0_196 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c196
*+ bl_0_196 br_0_196 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c196
*+ bl_0_196 br_0_196 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c196
*+ bl_0_196 br_0_196 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c196
*+ bl_0_196 br_0_196 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c196
*+ bl_0_196 br_0_196 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c196
*+ bl_0_196 br_0_196 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c196
*+ bl_0_196 br_0_196 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c196
*+ bl_0_196 br_0_196 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c196
*+ bl_0_196 br_0_196 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c196
*+ bl_0_196 br_0_196 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c196
*+ bl_0_196 br_0_196 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c196
*+ bl_0_196 br_0_196 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c196
*+ bl_0_196 br_0_196 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c196
*+ bl_0_196 br_0_196 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c196
*+ bl_0_196 br_0_196 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c196
*+ bl_0_196 br_0_196 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c196
*+ bl_0_196 br_0_196 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c196
*+ bl_0_196 br_0_196 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c196
*+ bl_0_196 br_0_196 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c196
*+ bl_0_196 br_0_196 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c196
*+ bl_0_196 br_0_196 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c196
*+ bl_0_196 br_0_196 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c196
*+ bl_0_196 br_0_196 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c196
*+ bl_0_196 br_0_196 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c196
*+ bl_0_196 br_0_196 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c196
*+ bl_0_196 br_0_196 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c196
*+ bl_0_196 br_0_196 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c196
*+ bl_0_196 br_0_196 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c196
*+ bl_0_196 br_0_196 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c196
*+ bl_0_196 br_0_196 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c196
*+ bl_0_196 br_0_196 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c196
*+ bl_0_196 br_0_196 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c196
*+ bl_0_196 br_0_196 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c196
*+ bl_0_196 br_0_196 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c196
*+ bl_0_196 br_0_196 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c196
+ bl_0_196 br_0_196 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c197
+ bl_0_197 br_0_197 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c197
*+ bl_0_197 br_0_197 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c197
*+ bl_0_197 br_0_197 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c197
*+ bl_0_197 br_0_197 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c197
*+ bl_0_197 br_0_197 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c197
*+ bl_0_197 br_0_197 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c197
*+ bl_0_197 br_0_197 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c197
*+ bl_0_197 br_0_197 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c197
*+ bl_0_197 br_0_197 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c197
*+ bl_0_197 br_0_197 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c197
*+ bl_0_197 br_0_197 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c197
*+ bl_0_197 br_0_197 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c197
*+ bl_0_197 br_0_197 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c197
*+ bl_0_197 br_0_197 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c197
*+ bl_0_197 br_0_197 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c197
*+ bl_0_197 br_0_197 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c197
*+ bl_0_197 br_0_197 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c197
*+ bl_0_197 br_0_197 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c197
*+ bl_0_197 br_0_197 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c197
*+ bl_0_197 br_0_197 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c197
*+ bl_0_197 br_0_197 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c197
*+ bl_0_197 br_0_197 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c197
*+ bl_0_197 br_0_197 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c197
*+ bl_0_197 br_0_197 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c197
*+ bl_0_197 br_0_197 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c197
*+ bl_0_197 br_0_197 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c197
*+ bl_0_197 br_0_197 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c197
*+ bl_0_197 br_0_197 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c197
*+ bl_0_197 br_0_197 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c197
*+ bl_0_197 br_0_197 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c197
*+ bl_0_197 br_0_197 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c197
*+ bl_0_197 br_0_197 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c197
*+ bl_0_197 br_0_197 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c197
*+ bl_0_197 br_0_197 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c197
*+ bl_0_197 br_0_197 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c197
*+ bl_0_197 br_0_197 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c197
*+ bl_0_197 br_0_197 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c197
*+ bl_0_197 br_0_197 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c197
*+ bl_0_197 br_0_197 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c197
*+ bl_0_197 br_0_197 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c197
*+ bl_0_197 br_0_197 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c197
*+ bl_0_197 br_0_197 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c197
*+ bl_0_197 br_0_197 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c197
*+ bl_0_197 br_0_197 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c197
*+ bl_0_197 br_0_197 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c197
*+ bl_0_197 br_0_197 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c197
*+ bl_0_197 br_0_197 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c197
*+ bl_0_197 br_0_197 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c197
*+ bl_0_197 br_0_197 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c197
*+ bl_0_197 br_0_197 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c197
*+ bl_0_197 br_0_197 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c197
*+ bl_0_197 br_0_197 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c197
*+ bl_0_197 br_0_197 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c197
*+ bl_0_197 br_0_197 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c197
*+ bl_0_197 br_0_197 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c197
*+ bl_0_197 br_0_197 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c197
*+ bl_0_197 br_0_197 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c197
*+ bl_0_197 br_0_197 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c197
*+ bl_0_197 br_0_197 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c197
*+ bl_0_197 br_0_197 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c197
*+ bl_0_197 br_0_197 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c197
*+ bl_0_197 br_0_197 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c197
*+ bl_0_197 br_0_197 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c197
*+ bl_0_197 br_0_197 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c197
*+ bl_0_197 br_0_197 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c197
*+ bl_0_197 br_0_197 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c197
*+ bl_0_197 br_0_197 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c197
*+ bl_0_197 br_0_197 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c197
*+ bl_0_197 br_0_197 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c197
*+ bl_0_197 br_0_197 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c197
*+ bl_0_197 br_0_197 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c197
*+ bl_0_197 br_0_197 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c197
*+ bl_0_197 br_0_197 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c197
*+ bl_0_197 br_0_197 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c197
*+ bl_0_197 br_0_197 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c197
*+ bl_0_197 br_0_197 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c197
*+ bl_0_197 br_0_197 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c197
*+ bl_0_197 br_0_197 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c197
*+ bl_0_197 br_0_197 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c197
*+ bl_0_197 br_0_197 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c197
*+ bl_0_197 br_0_197 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c197
*+ bl_0_197 br_0_197 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c197
*+ bl_0_197 br_0_197 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c197
*+ bl_0_197 br_0_197 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c197
*+ bl_0_197 br_0_197 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c197
*+ bl_0_197 br_0_197 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c197
*+ bl_0_197 br_0_197 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c197
*+ bl_0_197 br_0_197 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c197
*+ bl_0_197 br_0_197 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c197
*+ bl_0_197 br_0_197 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c197
*+ bl_0_197 br_0_197 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c197
*+ bl_0_197 br_0_197 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c197
*+ bl_0_197 br_0_197 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c197
*+ bl_0_197 br_0_197 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c197
*+ bl_0_197 br_0_197 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c197
*+ bl_0_197 br_0_197 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c197
*+ bl_0_197 br_0_197 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c197
*+ bl_0_197 br_0_197 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c197
*+ bl_0_197 br_0_197 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c197
*+ bl_0_197 br_0_197 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c197
*+ bl_0_197 br_0_197 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c197
*+ bl_0_197 br_0_197 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c197
*+ bl_0_197 br_0_197 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c197
*+ bl_0_197 br_0_197 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c197
*+ bl_0_197 br_0_197 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c197
*+ bl_0_197 br_0_197 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c197
*+ bl_0_197 br_0_197 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c197
*+ bl_0_197 br_0_197 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c197
*+ bl_0_197 br_0_197 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c197
*+ bl_0_197 br_0_197 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c197
*+ bl_0_197 br_0_197 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c197
*+ bl_0_197 br_0_197 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c197
*+ bl_0_197 br_0_197 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c197
*+ bl_0_197 br_0_197 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c197
*+ bl_0_197 br_0_197 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c197
*+ bl_0_197 br_0_197 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c197
*+ bl_0_197 br_0_197 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c197
*+ bl_0_197 br_0_197 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c197
*+ bl_0_197 br_0_197 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c197
*+ bl_0_197 br_0_197 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c197
*+ bl_0_197 br_0_197 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c197
*+ bl_0_197 br_0_197 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c197
*+ bl_0_197 br_0_197 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c197
*+ bl_0_197 br_0_197 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c197
*+ bl_0_197 br_0_197 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c197
*+ bl_0_197 br_0_197 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c197
*+ bl_0_197 br_0_197 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c197
+ bl_0_197 br_0_197 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c198
+ bl_0_198 br_0_198 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c198
*+ bl_0_198 br_0_198 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c198
*+ bl_0_198 br_0_198 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c198
*+ bl_0_198 br_0_198 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c198
*+ bl_0_198 br_0_198 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c198
*+ bl_0_198 br_0_198 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c198
*+ bl_0_198 br_0_198 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c198
*+ bl_0_198 br_0_198 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c198
*+ bl_0_198 br_0_198 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c198
*+ bl_0_198 br_0_198 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c198
*+ bl_0_198 br_0_198 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c198
*+ bl_0_198 br_0_198 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c198
*+ bl_0_198 br_0_198 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c198
*+ bl_0_198 br_0_198 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c198
*+ bl_0_198 br_0_198 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c198
*+ bl_0_198 br_0_198 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c198
*+ bl_0_198 br_0_198 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c198
*+ bl_0_198 br_0_198 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c198
*+ bl_0_198 br_0_198 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c198
*+ bl_0_198 br_0_198 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c198
*+ bl_0_198 br_0_198 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c198
*+ bl_0_198 br_0_198 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c198
*+ bl_0_198 br_0_198 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c198
*+ bl_0_198 br_0_198 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c198
*+ bl_0_198 br_0_198 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c198
*+ bl_0_198 br_0_198 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c198
*+ bl_0_198 br_0_198 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c198
*+ bl_0_198 br_0_198 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c198
*+ bl_0_198 br_0_198 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c198
*+ bl_0_198 br_0_198 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c198
*+ bl_0_198 br_0_198 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c198
*+ bl_0_198 br_0_198 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c198
*+ bl_0_198 br_0_198 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c198
*+ bl_0_198 br_0_198 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c198
*+ bl_0_198 br_0_198 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c198
*+ bl_0_198 br_0_198 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c198
*+ bl_0_198 br_0_198 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c198
*+ bl_0_198 br_0_198 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c198
*+ bl_0_198 br_0_198 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c198
*+ bl_0_198 br_0_198 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c198
*+ bl_0_198 br_0_198 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c198
*+ bl_0_198 br_0_198 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c198
*+ bl_0_198 br_0_198 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c198
*+ bl_0_198 br_0_198 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c198
*+ bl_0_198 br_0_198 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c198
*+ bl_0_198 br_0_198 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c198
*+ bl_0_198 br_0_198 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c198
*+ bl_0_198 br_0_198 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c198
*+ bl_0_198 br_0_198 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c198
*+ bl_0_198 br_0_198 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c198
*+ bl_0_198 br_0_198 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c198
*+ bl_0_198 br_0_198 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c198
*+ bl_0_198 br_0_198 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c198
*+ bl_0_198 br_0_198 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c198
*+ bl_0_198 br_0_198 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c198
*+ bl_0_198 br_0_198 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c198
*+ bl_0_198 br_0_198 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c198
*+ bl_0_198 br_0_198 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c198
*+ bl_0_198 br_0_198 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c198
*+ bl_0_198 br_0_198 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c198
*+ bl_0_198 br_0_198 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c198
*+ bl_0_198 br_0_198 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c198
*+ bl_0_198 br_0_198 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c198
*+ bl_0_198 br_0_198 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c198
*+ bl_0_198 br_0_198 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c198
*+ bl_0_198 br_0_198 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c198
*+ bl_0_198 br_0_198 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c198
*+ bl_0_198 br_0_198 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c198
*+ bl_0_198 br_0_198 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c198
*+ bl_0_198 br_0_198 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c198
*+ bl_0_198 br_0_198 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c198
*+ bl_0_198 br_0_198 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c198
*+ bl_0_198 br_0_198 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c198
*+ bl_0_198 br_0_198 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c198
*+ bl_0_198 br_0_198 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c198
*+ bl_0_198 br_0_198 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c198
*+ bl_0_198 br_0_198 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c198
*+ bl_0_198 br_0_198 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c198
*+ bl_0_198 br_0_198 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c198
*+ bl_0_198 br_0_198 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c198
*+ bl_0_198 br_0_198 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c198
*+ bl_0_198 br_0_198 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c198
*+ bl_0_198 br_0_198 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c198
*+ bl_0_198 br_0_198 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c198
*+ bl_0_198 br_0_198 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c198
*+ bl_0_198 br_0_198 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c198
*+ bl_0_198 br_0_198 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c198
*+ bl_0_198 br_0_198 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c198
*+ bl_0_198 br_0_198 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c198
*+ bl_0_198 br_0_198 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c198
*+ bl_0_198 br_0_198 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c198
*+ bl_0_198 br_0_198 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c198
*+ bl_0_198 br_0_198 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c198
*+ bl_0_198 br_0_198 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c198
*+ bl_0_198 br_0_198 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c198
*+ bl_0_198 br_0_198 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c198
*+ bl_0_198 br_0_198 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c198
*+ bl_0_198 br_0_198 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c198
*+ bl_0_198 br_0_198 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c198
*+ bl_0_198 br_0_198 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c198
*+ bl_0_198 br_0_198 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c198
*+ bl_0_198 br_0_198 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c198
*+ bl_0_198 br_0_198 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c198
*+ bl_0_198 br_0_198 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c198
*+ bl_0_198 br_0_198 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c198
*+ bl_0_198 br_0_198 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c198
*+ bl_0_198 br_0_198 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c198
*+ bl_0_198 br_0_198 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c198
*+ bl_0_198 br_0_198 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c198
*+ bl_0_198 br_0_198 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c198
*+ bl_0_198 br_0_198 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c198
*+ bl_0_198 br_0_198 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c198
*+ bl_0_198 br_0_198 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c198
*+ bl_0_198 br_0_198 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c198
*+ bl_0_198 br_0_198 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c198
*+ bl_0_198 br_0_198 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c198
*+ bl_0_198 br_0_198 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c198
*+ bl_0_198 br_0_198 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c198
*+ bl_0_198 br_0_198 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c198
*+ bl_0_198 br_0_198 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c198
*+ bl_0_198 br_0_198 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c198
*+ bl_0_198 br_0_198 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c198
*+ bl_0_198 br_0_198 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c198
*+ bl_0_198 br_0_198 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c198
*+ bl_0_198 br_0_198 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c198
*+ bl_0_198 br_0_198 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c198
*+ bl_0_198 br_0_198 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c198
+ bl_0_198 br_0_198 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c199
+ bl_0_199 br_0_199 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c199
*+ bl_0_199 br_0_199 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c199
*+ bl_0_199 br_0_199 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c199
*+ bl_0_199 br_0_199 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c199
*+ bl_0_199 br_0_199 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c199
*+ bl_0_199 br_0_199 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c199
*+ bl_0_199 br_0_199 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c199
*+ bl_0_199 br_0_199 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c199
*+ bl_0_199 br_0_199 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c199
*+ bl_0_199 br_0_199 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c199
*+ bl_0_199 br_0_199 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c199
*+ bl_0_199 br_0_199 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c199
*+ bl_0_199 br_0_199 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c199
*+ bl_0_199 br_0_199 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c199
*+ bl_0_199 br_0_199 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c199
*+ bl_0_199 br_0_199 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c199
*+ bl_0_199 br_0_199 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c199
*+ bl_0_199 br_0_199 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c199
*+ bl_0_199 br_0_199 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c199
*+ bl_0_199 br_0_199 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c199
*+ bl_0_199 br_0_199 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c199
*+ bl_0_199 br_0_199 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c199
*+ bl_0_199 br_0_199 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c199
*+ bl_0_199 br_0_199 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c199
*+ bl_0_199 br_0_199 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c199
*+ bl_0_199 br_0_199 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c199
*+ bl_0_199 br_0_199 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c199
*+ bl_0_199 br_0_199 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c199
*+ bl_0_199 br_0_199 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c199
*+ bl_0_199 br_0_199 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c199
*+ bl_0_199 br_0_199 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c199
*+ bl_0_199 br_0_199 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c199
*+ bl_0_199 br_0_199 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c199
*+ bl_0_199 br_0_199 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c199
*+ bl_0_199 br_0_199 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c199
*+ bl_0_199 br_0_199 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c199
*+ bl_0_199 br_0_199 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c199
*+ bl_0_199 br_0_199 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c199
*+ bl_0_199 br_0_199 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c199
*+ bl_0_199 br_0_199 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c199
*+ bl_0_199 br_0_199 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c199
*+ bl_0_199 br_0_199 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c199
*+ bl_0_199 br_0_199 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c199
*+ bl_0_199 br_0_199 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c199
*+ bl_0_199 br_0_199 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c199
*+ bl_0_199 br_0_199 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c199
*+ bl_0_199 br_0_199 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c199
*+ bl_0_199 br_0_199 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c199
*+ bl_0_199 br_0_199 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c199
*+ bl_0_199 br_0_199 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c199
*+ bl_0_199 br_0_199 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c199
*+ bl_0_199 br_0_199 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c199
*+ bl_0_199 br_0_199 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c199
*+ bl_0_199 br_0_199 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c199
*+ bl_0_199 br_0_199 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c199
*+ bl_0_199 br_0_199 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c199
*+ bl_0_199 br_0_199 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c199
*+ bl_0_199 br_0_199 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c199
*+ bl_0_199 br_0_199 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c199
*+ bl_0_199 br_0_199 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c199
*+ bl_0_199 br_0_199 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c199
*+ bl_0_199 br_0_199 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c199
*+ bl_0_199 br_0_199 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c199
*+ bl_0_199 br_0_199 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c199
*+ bl_0_199 br_0_199 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c199
*+ bl_0_199 br_0_199 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c199
*+ bl_0_199 br_0_199 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c199
*+ bl_0_199 br_0_199 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c199
*+ bl_0_199 br_0_199 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c199
*+ bl_0_199 br_0_199 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c199
*+ bl_0_199 br_0_199 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c199
*+ bl_0_199 br_0_199 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c199
*+ bl_0_199 br_0_199 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c199
*+ bl_0_199 br_0_199 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c199
*+ bl_0_199 br_0_199 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c199
*+ bl_0_199 br_0_199 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c199
*+ bl_0_199 br_0_199 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c199
*+ bl_0_199 br_0_199 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c199
*+ bl_0_199 br_0_199 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c199
*+ bl_0_199 br_0_199 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c199
*+ bl_0_199 br_0_199 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c199
*+ bl_0_199 br_0_199 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c199
*+ bl_0_199 br_0_199 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c199
*+ bl_0_199 br_0_199 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c199
*+ bl_0_199 br_0_199 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c199
*+ bl_0_199 br_0_199 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c199
*+ bl_0_199 br_0_199 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c199
*+ bl_0_199 br_0_199 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c199
*+ bl_0_199 br_0_199 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c199
*+ bl_0_199 br_0_199 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c199
*+ bl_0_199 br_0_199 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c199
*+ bl_0_199 br_0_199 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c199
*+ bl_0_199 br_0_199 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c199
*+ bl_0_199 br_0_199 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c199
*+ bl_0_199 br_0_199 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c199
*+ bl_0_199 br_0_199 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c199
*+ bl_0_199 br_0_199 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c199
*+ bl_0_199 br_0_199 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c199
*+ bl_0_199 br_0_199 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c199
*+ bl_0_199 br_0_199 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c199
*+ bl_0_199 br_0_199 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c199
*+ bl_0_199 br_0_199 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c199
*+ bl_0_199 br_0_199 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c199
*+ bl_0_199 br_0_199 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c199
*+ bl_0_199 br_0_199 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c199
*+ bl_0_199 br_0_199 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c199
*+ bl_0_199 br_0_199 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c199
*+ bl_0_199 br_0_199 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c199
*+ bl_0_199 br_0_199 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c199
*+ bl_0_199 br_0_199 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c199
*+ bl_0_199 br_0_199 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c199
*+ bl_0_199 br_0_199 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c199
*+ bl_0_199 br_0_199 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c199
*+ bl_0_199 br_0_199 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c199
*+ bl_0_199 br_0_199 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c199
*+ bl_0_199 br_0_199 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c199
*+ bl_0_199 br_0_199 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c199
*+ bl_0_199 br_0_199 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c199
*+ bl_0_199 br_0_199 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c199
*+ bl_0_199 br_0_199 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c199
*+ bl_0_199 br_0_199 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c199
*+ bl_0_199 br_0_199 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c199
*+ bl_0_199 br_0_199 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c199
*+ bl_0_199 br_0_199 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c199
*+ bl_0_199 br_0_199 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c199
*+ bl_0_199 br_0_199 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c199
*+ bl_0_199 br_0_199 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c199
+ bl_0_199 br_0_199 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c200
+ bl_0_200 br_0_200 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c200
*+ bl_0_200 br_0_200 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c200
*+ bl_0_200 br_0_200 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c200
*+ bl_0_200 br_0_200 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c200
*+ bl_0_200 br_0_200 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c200
*+ bl_0_200 br_0_200 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c200
*+ bl_0_200 br_0_200 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c200
*+ bl_0_200 br_0_200 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c200
*+ bl_0_200 br_0_200 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c200
*+ bl_0_200 br_0_200 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c200
*+ bl_0_200 br_0_200 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c200
*+ bl_0_200 br_0_200 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c200
*+ bl_0_200 br_0_200 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c200
*+ bl_0_200 br_0_200 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c200
*+ bl_0_200 br_0_200 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c200
*+ bl_0_200 br_0_200 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c200
*+ bl_0_200 br_0_200 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c200
*+ bl_0_200 br_0_200 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c200
*+ bl_0_200 br_0_200 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c200
*+ bl_0_200 br_0_200 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c200
*+ bl_0_200 br_0_200 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c200
*+ bl_0_200 br_0_200 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c200
*+ bl_0_200 br_0_200 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c200
*+ bl_0_200 br_0_200 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c200
*+ bl_0_200 br_0_200 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c200
*+ bl_0_200 br_0_200 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c200
*+ bl_0_200 br_0_200 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c200
*+ bl_0_200 br_0_200 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c200
*+ bl_0_200 br_0_200 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c200
*+ bl_0_200 br_0_200 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c200
*+ bl_0_200 br_0_200 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c200
*+ bl_0_200 br_0_200 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c200
*+ bl_0_200 br_0_200 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c200
*+ bl_0_200 br_0_200 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c200
*+ bl_0_200 br_0_200 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c200
*+ bl_0_200 br_0_200 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c200
*+ bl_0_200 br_0_200 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c200
*+ bl_0_200 br_0_200 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c200
*+ bl_0_200 br_0_200 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c200
*+ bl_0_200 br_0_200 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c200
*+ bl_0_200 br_0_200 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c200
*+ bl_0_200 br_0_200 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c200
*+ bl_0_200 br_0_200 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c200
*+ bl_0_200 br_0_200 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c200
*+ bl_0_200 br_0_200 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c200
*+ bl_0_200 br_0_200 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c200
*+ bl_0_200 br_0_200 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c200
*+ bl_0_200 br_0_200 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c200
*+ bl_0_200 br_0_200 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c200
*+ bl_0_200 br_0_200 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c200
*+ bl_0_200 br_0_200 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c200
*+ bl_0_200 br_0_200 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c200
*+ bl_0_200 br_0_200 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c200
*+ bl_0_200 br_0_200 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c200
*+ bl_0_200 br_0_200 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c200
*+ bl_0_200 br_0_200 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c200
*+ bl_0_200 br_0_200 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c200
*+ bl_0_200 br_0_200 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c200
*+ bl_0_200 br_0_200 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c200
*+ bl_0_200 br_0_200 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c200
*+ bl_0_200 br_0_200 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c200
*+ bl_0_200 br_0_200 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c200
*+ bl_0_200 br_0_200 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c200
*+ bl_0_200 br_0_200 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c200
*+ bl_0_200 br_0_200 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c200
*+ bl_0_200 br_0_200 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c200
*+ bl_0_200 br_0_200 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c200
*+ bl_0_200 br_0_200 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c200
*+ bl_0_200 br_0_200 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c200
*+ bl_0_200 br_0_200 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c200
*+ bl_0_200 br_0_200 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c200
*+ bl_0_200 br_0_200 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c200
*+ bl_0_200 br_0_200 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c200
*+ bl_0_200 br_0_200 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c200
*+ bl_0_200 br_0_200 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c200
*+ bl_0_200 br_0_200 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c200
*+ bl_0_200 br_0_200 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c200
*+ bl_0_200 br_0_200 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c200
*+ bl_0_200 br_0_200 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c200
*+ bl_0_200 br_0_200 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c200
*+ bl_0_200 br_0_200 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c200
*+ bl_0_200 br_0_200 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c200
*+ bl_0_200 br_0_200 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c200
*+ bl_0_200 br_0_200 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c200
*+ bl_0_200 br_0_200 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c200
*+ bl_0_200 br_0_200 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c200
*+ bl_0_200 br_0_200 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c200
*+ bl_0_200 br_0_200 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c200
*+ bl_0_200 br_0_200 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c200
*+ bl_0_200 br_0_200 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c200
*+ bl_0_200 br_0_200 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c200
*+ bl_0_200 br_0_200 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c200
*+ bl_0_200 br_0_200 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c200
*+ bl_0_200 br_0_200 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c200
*+ bl_0_200 br_0_200 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c200
*+ bl_0_200 br_0_200 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c200
*+ bl_0_200 br_0_200 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c200
*+ bl_0_200 br_0_200 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c200
*+ bl_0_200 br_0_200 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c200
*+ bl_0_200 br_0_200 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c200
*+ bl_0_200 br_0_200 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c200
*+ bl_0_200 br_0_200 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c200
*+ bl_0_200 br_0_200 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c200
*+ bl_0_200 br_0_200 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c200
*+ bl_0_200 br_0_200 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c200
*+ bl_0_200 br_0_200 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c200
*+ bl_0_200 br_0_200 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c200
*+ bl_0_200 br_0_200 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c200
*+ bl_0_200 br_0_200 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c200
*+ bl_0_200 br_0_200 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c200
*+ bl_0_200 br_0_200 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c200
*+ bl_0_200 br_0_200 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c200
*+ bl_0_200 br_0_200 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c200
*+ bl_0_200 br_0_200 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c200
*+ bl_0_200 br_0_200 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c200
*+ bl_0_200 br_0_200 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c200
*+ bl_0_200 br_0_200 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c200
*+ bl_0_200 br_0_200 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c200
*+ bl_0_200 br_0_200 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c200
*+ bl_0_200 br_0_200 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c200
*+ bl_0_200 br_0_200 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c200
*+ bl_0_200 br_0_200 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c200
*+ bl_0_200 br_0_200 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c200
*+ bl_0_200 br_0_200 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c200
*+ bl_0_200 br_0_200 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c200
*+ bl_0_200 br_0_200 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c200
*+ bl_0_200 br_0_200 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c200
+ bl_0_200 br_0_200 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c201
+ bl_0_201 br_0_201 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c201
*+ bl_0_201 br_0_201 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c201
*+ bl_0_201 br_0_201 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c201
*+ bl_0_201 br_0_201 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c201
*+ bl_0_201 br_0_201 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c201
*+ bl_0_201 br_0_201 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c201
*+ bl_0_201 br_0_201 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c201
*+ bl_0_201 br_0_201 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c201
*+ bl_0_201 br_0_201 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c201
*+ bl_0_201 br_0_201 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c201
*+ bl_0_201 br_0_201 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c201
*+ bl_0_201 br_0_201 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c201
*+ bl_0_201 br_0_201 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c201
*+ bl_0_201 br_0_201 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c201
*+ bl_0_201 br_0_201 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c201
*+ bl_0_201 br_0_201 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c201
*+ bl_0_201 br_0_201 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c201
*+ bl_0_201 br_0_201 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c201
*+ bl_0_201 br_0_201 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c201
*+ bl_0_201 br_0_201 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c201
*+ bl_0_201 br_0_201 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c201
*+ bl_0_201 br_0_201 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c201
*+ bl_0_201 br_0_201 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c201
*+ bl_0_201 br_0_201 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c201
*+ bl_0_201 br_0_201 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c201
*+ bl_0_201 br_0_201 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c201
*+ bl_0_201 br_0_201 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c201
*+ bl_0_201 br_0_201 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c201
*+ bl_0_201 br_0_201 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c201
*+ bl_0_201 br_0_201 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c201
*+ bl_0_201 br_0_201 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c201
*+ bl_0_201 br_0_201 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c201
*+ bl_0_201 br_0_201 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c201
*+ bl_0_201 br_0_201 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c201
*+ bl_0_201 br_0_201 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c201
*+ bl_0_201 br_0_201 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c201
*+ bl_0_201 br_0_201 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c201
*+ bl_0_201 br_0_201 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c201
*+ bl_0_201 br_0_201 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c201
*+ bl_0_201 br_0_201 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c201
*+ bl_0_201 br_0_201 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c201
*+ bl_0_201 br_0_201 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c201
*+ bl_0_201 br_0_201 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c201
*+ bl_0_201 br_0_201 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c201
*+ bl_0_201 br_0_201 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c201
*+ bl_0_201 br_0_201 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c201
*+ bl_0_201 br_0_201 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c201
*+ bl_0_201 br_0_201 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c201
*+ bl_0_201 br_0_201 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c201
*+ bl_0_201 br_0_201 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c201
*+ bl_0_201 br_0_201 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c201
*+ bl_0_201 br_0_201 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c201
*+ bl_0_201 br_0_201 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c201
*+ bl_0_201 br_0_201 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c201
*+ bl_0_201 br_0_201 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c201
*+ bl_0_201 br_0_201 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c201
*+ bl_0_201 br_0_201 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c201
*+ bl_0_201 br_0_201 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c201
*+ bl_0_201 br_0_201 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c201
*+ bl_0_201 br_0_201 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c201
*+ bl_0_201 br_0_201 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c201
*+ bl_0_201 br_0_201 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c201
*+ bl_0_201 br_0_201 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c201
*+ bl_0_201 br_0_201 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c201
*+ bl_0_201 br_0_201 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c201
*+ bl_0_201 br_0_201 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c201
*+ bl_0_201 br_0_201 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c201
*+ bl_0_201 br_0_201 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c201
*+ bl_0_201 br_0_201 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c201
*+ bl_0_201 br_0_201 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c201
*+ bl_0_201 br_0_201 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c201
*+ bl_0_201 br_0_201 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c201
*+ bl_0_201 br_0_201 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c201
*+ bl_0_201 br_0_201 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c201
*+ bl_0_201 br_0_201 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c201
*+ bl_0_201 br_0_201 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c201
*+ bl_0_201 br_0_201 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c201
*+ bl_0_201 br_0_201 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c201
*+ bl_0_201 br_0_201 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c201
*+ bl_0_201 br_0_201 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c201
*+ bl_0_201 br_0_201 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c201
*+ bl_0_201 br_0_201 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c201
*+ bl_0_201 br_0_201 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c201
*+ bl_0_201 br_0_201 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c201
*+ bl_0_201 br_0_201 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c201
*+ bl_0_201 br_0_201 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c201
*+ bl_0_201 br_0_201 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c201
*+ bl_0_201 br_0_201 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c201
*+ bl_0_201 br_0_201 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c201
*+ bl_0_201 br_0_201 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c201
*+ bl_0_201 br_0_201 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c201
*+ bl_0_201 br_0_201 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c201
*+ bl_0_201 br_0_201 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c201
*+ bl_0_201 br_0_201 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c201
*+ bl_0_201 br_0_201 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c201
*+ bl_0_201 br_0_201 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c201
*+ bl_0_201 br_0_201 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c201
*+ bl_0_201 br_0_201 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c201
*+ bl_0_201 br_0_201 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c201
*+ bl_0_201 br_0_201 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c201
*+ bl_0_201 br_0_201 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c201
*+ bl_0_201 br_0_201 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c201
*+ bl_0_201 br_0_201 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c201
*+ bl_0_201 br_0_201 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c201
*+ bl_0_201 br_0_201 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c201
*+ bl_0_201 br_0_201 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c201
*+ bl_0_201 br_0_201 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c201
*+ bl_0_201 br_0_201 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c201
*+ bl_0_201 br_0_201 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c201
*+ bl_0_201 br_0_201 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c201
*+ bl_0_201 br_0_201 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c201
*+ bl_0_201 br_0_201 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c201
*+ bl_0_201 br_0_201 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c201
*+ bl_0_201 br_0_201 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c201
*+ bl_0_201 br_0_201 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c201
*+ bl_0_201 br_0_201 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c201
*+ bl_0_201 br_0_201 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c201
*+ bl_0_201 br_0_201 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c201
*+ bl_0_201 br_0_201 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c201
*+ bl_0_201 br_0_201 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c201
*+ bl_0_201 br_0_201 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c201
*+ bl_0_201 br_0_201 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c201
*+ bl_0_201 br_0_201 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c201
*+ bl_0_201 br_0_201 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c201
*+ bl_0_201 br_0_201 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c201
*+ bl_0_201 br_0_201 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c201
*+ bl_0_201 br_0_201 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c201
+ bl_0_201 br_0_201 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c202
+ bl_0_202 br_0_202 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c202
*+ bl_0_202 br_0_202 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c202
*+ bl_0_202 br_0_202 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c202
*+ bl_0_202 br_0_202 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c202
*+ bl_0_202 br_0_202 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c202
*+ bl_0_202 br_0_202 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c202
*+ bl_0_202 br_0_202 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c202
*+ bl_0_202 br_0_202 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c202
*+ bl_0_202 br_0_202 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c202
*+ bl_0_202 br_0_202 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c202
*+ bl_0_202 br_0_202 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c202
*+ bl_0_202 br_0_202 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c202
*+ bl_0_202 br_0_202 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c202
*+ bl_0_202 br_0_202 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c202
*+ bl_0_202 br_0_202 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c202
*+ bl_0_202 br_0_202 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c202
*+ bl_0_202 br_0_202 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c202
*+ bl_0_202 br_0_202 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c202
*+ bl_0_202 br_0_202 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c202
*+ bl_0_202 br_0_202 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c202
*+ bl_0_202 br_0_202 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c202
*+ bl_0_202 br_0_202 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c202
*+ bl_0_202 br_0_202 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c202
*+ bl_0_202 br_0_202 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c202
*+ bl_0_202 br_0_202 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c202
*+ bl_0_202 br_0_202 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c202
*+ bl_0_202 br_0_202 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c202
*+ bl_0_202 br_0_202 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c202
*+ bl_0_202 br_0_202 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c202
*+ bl_0_202 br_0_202 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c202
*+ bl_0_202 br_0_202 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c202
*+ bl_0_202 br_0_202 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c202
*+ bl_0_202 br_0_202 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c202
*+ bl_0_202 br_0_202 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c202
*+ bl_0_202 br_0_202 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c202
*+ bl_0_202 br_0_202 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c202
*+ bl_0_202 br_0_202 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c202
*+ bl_0_202 br_0_202 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c202
*+ bl_0_202 br_0_202 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c202
*+ bl_0_202 br_0_202 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c202
*+ bl_0_202 br_0_202 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c202
*+ bl_0_202 br_0_202 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c202
*+ bl_0_202 br_0_202 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c202
*+ bl_0_202 br_0_202 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c202
*+ bl_0_202 br_0_202 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c202
*+ bl_0_202 br_0_202 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c202
*+ bl_0_202 br_0_202 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c202
*+ bl_0_202 br_0_202 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c202
*+ bl_0_202 br_0_202 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c202
*+ bl_0_202 br_0_202 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c202
*+ bl_0_202 br_0_202 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c202
*+ bl_0_202 br_0_202 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c202
*+ bl_0_202 br_0_202 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c202
*+ bl_0_202 br_0_202 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c202
*+ bl_0_202 br_0_202 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c202
*+ bl_0_202 br_0_202 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c202
*+ bl_0_202 br_0_202 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c202
*+ bl_0_202 br_0_202 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c202
*+ bl_0_202 br_0_202 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c202
*+ bl_0_202 br_0_202 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c202
*+ bl_0_202 br_0_202 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c202
*+ bl_0_202 br_0_202 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c202
*+ bl_0_202 br_0_202 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c202
*+ bl_0_202 br_0_202 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c202
*+ bl_0_202 br_0_202 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c202
*+ bl_0_202 br_0_202 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c202
*+ bl_0_202 br_0_202 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c202
*+ bl_0_202 br_0_202 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c202
*+ bl_0_202 br_0_202 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c202
*+ bl_0_202 br_0_202 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c202
*+ bl_0_202 br_0_202 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c202
*+ bl_0_202 br_0_202 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c202
*+ bl_0_202 br_0_202 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c202
*+ bl_0_202 br_0_202 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c202
*+ bl_0_202 br_0_202 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c202
*+ bl_0_202 br_0_202 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c202
*+ bl_0_202 br_0_202 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c202
*+ bl_0_202 br_0_202 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c202
*+ bl_0_202 br_0_202 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c202
*+ bl_0_202 br_0_202 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c202
*+ bl_0_202 br_0_202 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c202
*+ bl_0_202 br_0_202 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c202
*+ bl_0_202 br_0_202 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c202
*+ bl_0_202 br_0_202 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c202
*+ bl_0_202 br_0_202 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c202
*+ bl_0_202 br_0_202 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c202
*+ bl_0_202 br_0_202 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c202
*+ bl_0_202 br_0_202 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c202
*+ bl_0_202 br_0_202 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c202
*+ bl_0_202 br_0_202 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c202
*+ bl_0_202 br_0_202 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c202
*+ bl_0_202 br_0_202 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c202
*+ bl_0_202 br_0_202 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c202
*+ bl_0_202 br_0_202 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c202
*+ bl_0_202 br_0_202 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c202
*+ bl_0_202 br_0_202 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c202
*+ bl_0_202 br_0_202 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c202
*+ bl_0_202 br_0_202 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c202
*+ bl_0_202 br_0_202 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c202
*+ bl_0_202 br_0_202 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c202
*+ bl_0_202 br_0_202 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c202
*+ bl_0_202 br_0_202 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c202
*+ bl_0_202 br_0_202 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c202
*+ bl_0_202 br_0_202 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c202
*+ bl_0_202 br_0_202 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c202
*+ bl_0_202 br_0_202 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c202
*+ bl_0_202 br_0_202 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c202
*+ bl_0_202 br_0_202 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c202
*+ bl_0_202 br_0_202 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c202
*+ bl_0_202 br_0_202 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c202
*+ bl_0_202 br_0_202 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c202
*+ bl_0_202 br_0_202 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c202
*+ bl_0_202 br_0_202 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c202
*+ bl_0_202 br_0_202 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c202
*+ bl_0_202 br_0_202 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c202
*+ bl_0_202 br_0_202 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c202
*+ bl_0_202 br_0_202 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c202
*+ bl_0_202 br_0_202 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c202
*+ bl_0_202 br_0_202 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c202
*+ bl_0_202 br_0_202 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c202
*+ bl_0_202 br_0_202 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c202
*+ bl_0_202 br_0_202 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c202
*+ bl_0_202 br_0_202 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c202
*+ bl_0_202 br_0_202 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c202
*+ bl_0_202 br_0_202 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c202
*+ bl_0_202 br_0_202 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c202
*+ bl_0_202 br_0_202 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c202
+ bl_0_202 br_0_202 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c203
+ bl_0_203 br_0_203 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c203
*+ bl_0_203 br_0_203 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c203
*+ bl_0_203 br_0_203 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c203
*+ bl_0_203 br_0_203 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c203
*+ bl_0_203 br_0_203 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c203
*+ bl_0_203 br_0_203 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c203
*+ bl_0_203 br_0_203 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c203
*+ bl_0_203 br_0_203 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c203
*+ bl_0_203 br_0_203 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c203
*+ bl_0_203 br_0_203 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c203
*+ bl_0_203 br_0_203 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c203
*+ bl_0_203 br_0_203 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c203
*+ bl_0_203 br_0_203 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c203
*+ bl_0_203 br_0_203 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c203
*+ bl_0_203 br_0_203 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c203
*+ bl_0_203 br_0_203 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c203
*+ bl_0_203 br_0_203 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c203
*+ bl_0_203 br_0_203 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c203
*+ bl_0_203 br_0_203 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c203
*+ bl_0_203 br_0_203 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c203
*+ bl_0_203 br_0_203 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c203
*+ bl_0_203 br_0_203 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c203
*+ bl_0_203 br_0_203 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c203
*+ bl_0_203 br_0_203 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c203
*+ bl_0_203 br_0_203 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c203
*+ bl_0_203 br_0_203 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c203
*+ bl_0_203 br_0_203 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c203
*+ bl_0_203 br_0_203 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c203
*+ bl_0_203 br_0_203 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c203
*+ bl_0_203 br_0_203 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c203
*+ bl_0_203 br_0_203 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c203
*+ bl_0_203 br_0_203 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c203
*+ bl_0_203 br_0_203 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c203
*+ bl_0_203 br_0_203 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c203
*+ bl_0_203 br_0_203 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c203
*+ bl_0_203 br_0_203 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c203
*+ bl_0_203 br_0_203 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c203
*+ bl_0_203 br_0_203 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c203
*+ bl_0_203 br_0_203 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c203
*+ bl_0_203 br_0_203 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c203
*+ bl_0_203 br_0_203 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c203
*+ bl_0_203 br_0_203 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c203
*+ bl_0_203 br_0_203 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c203
*+ bl_0_203 br_0_203 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c203
*+ bl_0_203 br_0_203 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c203
*+ bl_0_203 br_0_203 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c203
*+ bl_0_203 br_0_203 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c203
*+ bl_0_203 br_0_203 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c203
*+ bl_0_203 br_0_203 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c203
*+ bl_0_203 br_0_203 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c203
*+ bl_0_203 br_0_203 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c203
*+ bl_0_203 br_0_203 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c203
*+ bl_0_203 br_0_203 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c203
*+ bl_0_203 br_0_203 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c203
*+ bl_0_203 br_0_203 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c203
*+ bl_0_203 br_0_203 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c203
*+ bl_0_203 br_0_203 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c203
*+ bl_0_203 br_0_203 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c203
*+ bl_0_203 br_0_203 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c203
*+ bl_0_203 br_0_203 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c203
*+ bl_0_203 br_0_203 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c203
*+ bl_0_203 br_0_203 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c203
*+ bl_0_203 br_0_203 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c203
*+ bl_0_203 br_0_203 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c203
*+ bl_0_203 br_0_203 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c203
*+ bl_0_203 br_0_203 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c203
*+ bl_0_203 br_0_203 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c203
*+ bl_0_203 br_0_203 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c203
*+ bl_0_203 br_0_203 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c203
*+ bl_0_203 br_0_203 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c203
*+ bl_0_203 br_0_203 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c203
*+ bl_0_203 br_0_203 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c203
*+ bl_0_203 br_0_203 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c203
*+ bl_0_203 br_0_203 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c203
*+ bl_0_203 br_0_203 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c203
*+ bl_0_203 br_0_203 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c203
*+ bl_0_203 br_0_203 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c203
*+ bl_0_203 br_0_203 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c203
*+ bl_0_203 br_0_203 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c203
*+ bl_0_203 br_0_203 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c203
*+ bl_0_203 br_0_203 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c203
*+ bl_0_203 br_0_203 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c203
*+ bl_0_203 br_0_203 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c203
*+ bl_0_203 br_0_203 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c203
*+ bl_0_203 br_0_203 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c203
*+ bl_0_203 br_0_203 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c203
*+ bl_0_203 br_0_203 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c203
*+ bl_0_203 br_0_203 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c203
*+ bl_0_203 br_0_203 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c203
*+ bl_0_203 br_0_203 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c203
*+ bl_0_203 br_0_203 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c203
*+ bl_0_203 br_0_203 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c203
*+ bl_0_203 br_0_203 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c203
*+ bl_0_203 br_0_203 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c203
*+ bl_0_203 br_0_203 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c203
*+ bl_0_203 br_0_203 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c203
*+ bl_0_203 br_0_203 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c203
*+ bl_0_203 br_0_203 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c203
*+ bl_0_203 br_0_203 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c203
*+ bl_0_203 br_0_203 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c203
*+ bl_0_203 br_0_203 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c203
*+ bl_0_203 br_0_203 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c203
*+ bl_0_203 br_0_203 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c203
*+ bl_0_203 br_0_203 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c203
*+ bl_0_203 br_0_203 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c203
*+ bl_0_203 br_0_203 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c203
*+ bl_0_203 br_0_203 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c203
*+ bl_0_203 br_0_203 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c203
*+ bl_0_203 br_0_203 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c203
*+ bl_0_203 br_0_203 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c203
*+ bl_0_203 br_0_203 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c203
*+ bl_0_203 br_0_203 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c203
*+ bl_0_203 br_0_203 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c203
*+ bl_0_203 br_0_203 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c203
*+ bl_0_203 br_0_203 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c203
*+ bl_0_203 br_0_203 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c203
*+ bl_0_203 br_0_203 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c203
*+ bl_0_203 br_0_203 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c203
*+ bl_0_203 br_0_203 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c203
*+ bl_0_203 br_0_203 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c203
*+ bl_0_203 br_0_203 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c203
*+ bl_0_203 br_0_203 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c203
*+ bl_0_203 br_0_203 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c203
*+ bl_0_203 br_0_203 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c203
*+ bl_0_203 br_0_203 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c203
*+ bl_0_203 br_0_203 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c203
*+ bl_0_203 br_0_203 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c203
+ bl_0_203 br_0_203 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c204
+ bl_0_204 br_0_204 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c204
*+ bl_0_204 br_0_204 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c204
*+ bl_0_204 br_0_204 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c204
*+ bl_0_204 br_0_204 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c204
*+ bl_0_204 br_0_204 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c204
*+ bl_0_204 br_0_204 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c204
*+ bl_0_204 br_0_204 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c204
*+ bl_0_204 br_0_204 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c204
*+ bl_0_204 br_0_204 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c204
*+ bl_0_204 br_0_204 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c204
*+ bl_0_204 br_0_204 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c204
*+ bl_0_204 br_0_204 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c204
*+ bl_0_204 br_0_204 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c204
*+ bl_0_204 br_0_204 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c204
*+ bl_0_204 br_0_204 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c204
*+ bl_0_204 br_0_204 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c204
*+ bl_0_204 br_0_204 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c204
*+ bl_0_204 br_0_204 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c204
*+ bl_0_204 br_0_204 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c204
*+ bl_0_204 br_0_204 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c204
*+ bl_0_204 br_0_204 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c204
*+ bl_0_204 br_0_204 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c204
*+ bl_0_204 br_0_204 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c204
*+ bl_0_204 br_0_204 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c204
*+ bl_0_204 br_0_204 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c204
*+ bl_0_204 br_0_204 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c204
*+ bl_0_204 br_0_204 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c204
*+ bl_0_204 br_0_204 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c204
*+ bl_0_204 br_0_204 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c204
*+ bl_0_204 br_0_204 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c204
*+ bl_0_204 br_0_204 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c204
*+ bl_0_204 br_0_204 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c204
*+ bl_0_204 br_0_204 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c204
*+ bl_0_204 br_0_204 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c204
*+ bl_0_204 br_0_204 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c204
*+ bl_0_204 br_0_204 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c204
*+ bl_0_204 br_0_204 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c204
*+ bl_0_204 br_0_204 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c204
*+ bl_0_204 br_0_204 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c204
*+ bl_0_204 br_0_204 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c204
*+ bl_0_204 br_0_204 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c204
*+ bl_0_204 br_0_204 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c204
*+ bl_0_204 br_0_204 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c204
*+ bl_0_204 br_0_204 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c204
*+ bl_0_204 br_0_204 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c204
*+ bl_0_204 br_0_204 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c204
*+ bl_0_204 br_0_204 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c204
*+ bl_0_204 br_0_204 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c204
*+ bl_0_204 br_0_204 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c204
*+ bl_0_204 br_0_204 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c204
*+ bl_0_204 br_0_204 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c204
*+ bl_0_204 br_0_204 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c204
*+ bl_0_204 br_0_204 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c204
*+ bl_0_204 br_0_204 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c204
*+ bl_0_204 br_0_204 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c204
*+ bl_0_204 br_0_204 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c204
*+ bl_0_204 br_0_204 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c204
*+ bl_0_204 br_0_204 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c204
*+ bl_0_204 br_0_204 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c204
*+ bl_0_204 br_0_204 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c204
*+ bl_0_204 br_0_204 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c204
*+ bl_0_204 br_0_204 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c204
*+ bl_0_204 br_0_204 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c204
*+ bl_0_204 br_0_204 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c204
*+ bl_0_204 br_0_204 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c204
*+ bl_0_204 br_0_204 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c204
*+ bl_0_204 br_0_204 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c204
*+ bl_0_204 br_0_204 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c204
*+ bl_0_204 br_0_204 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c204
*+ bl_0_204 br_0_204 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c204
*+ bl_0_204 br_0_204 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c204
*+ bl_0_204 br_0_204 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c204
*+ bl_0_204 br_0_204 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c204
*+ bl_0_204 br_0_204 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c204
*+ bl_0_204 br_0_204 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c204
*+ bl_0_204 br_0_204 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c204
*+ bl_0_204 br_0_204 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c204
*+ bl_0_204 br_0_204 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c204
*+ bl_0_204 br_0_204 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c204
*+ bl_0_204 br_0_204 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c204
*+ bl_0_204 br_0_204 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c204
*+ bl_0_204 br_0_204 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c204
*+ bl_0_204 br_0_204 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c204
*+ bl_0_204 br_0_204 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c204
*+ bl_0_204 br_0_204 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c204
*+ bl_0_204 br_0_204 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c204
*+ bl_0_204 br_0_204 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c204
*+ bl_0_204 br_0_204 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c204
*+ bl_0_204 br_0_204 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c204
*+ bl_0_204 br_0_204 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c204
*+ bl_0_204 br_0_204 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c204
*+ bl_0_204 br_0_204 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c204
*+ bl_0_204 br_0_204 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c204
*+ bl_0_204 br_0_204 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c204
*+ bl_0_204 br_0_204 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c204
*+ bl_0_204 br_0_204 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c204
*+ bl_0_204 br_0_204 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c204
*+ bl_0_204 br_0_204 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c204
*+ bl_0_204 br_0_204 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c204
*+ bl_0_204 br_0_204 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c204
*+ bl_0_204 br_0_204 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c204
*+ bl_0_204 br_0_204 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c204
*+ bl_0_204 br_0_204 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c204
*+ bl_0_204 br_0_204 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c204
*+ bl_0_204 br_0_204 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c204
*+ bl_0_204 br_0_204 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c204
*+ bl_0_204 br_0_204 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c204
*+ bl_0_204 br_0_204 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c204
*+ bl_0_204 br_0_204 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c204
*+ bl_0_204 br_0_204 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c204
*+ bl_0_204 br_0_204 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c204
*+ bl_0_204 br_0_204 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c204
*+ bl_0_204 br_0_204 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c204
*+ bl_0_204 br_0_204 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c204
*+ bl_0_204 br_0_204 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c204
*+ bl_0_204 br_0_204 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c204
*+ bl_0_204 br_0_204 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c204
*+ bl_0_204 br_0_204 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c204
*+ bl_0_204 br_0_204 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c204
*+ bl_0_204 br_0_204 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c204
*+ bl_0_204 br_0_204 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c204
*+ bl_0_204 br_0_204 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c204
*+ bl_0_204 br_0_204 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c204
*+ bl_0_204 br_0_204 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c204
*+ bl_0_204 br_0_204 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c204
*+ bl_0_204 br_0_204 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c204
*+ bl_0_204 br_0_204 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c204
+ bl_0_204 br_0_204 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c205
+ bl_0_205 br_0_205 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c205
*+ bl_0_205 br_0_205 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c205
*+ bl_0_205 br_0_205 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c205
*+ bl_0_205 br_0_205 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c205
*+ bl_0_205 br_0_205 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c205
*+ bl_0_205 br_0_205 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c205
*+ bl_0_205 br_0_205 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c205
*+ bl_0_205 br_0_205 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c205
*+ bl_0_205 br_0_205 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c205
*+ bl_0_205 br_0_205 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c205
*+ bl_0_205 br_0_205 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c205
*+ bl_0_205 br_0_205 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c205
*+ bl_0_205 br_0_205 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c205
*+ bl_0_205 br_0_205 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c205
*+ bl_0_205 br_0_205 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c205
*+ bl_0_205 br_0_205 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c205
*+ bl_0_205 br_0_205 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c205
*+ bl_0_205 br_0_205 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c205
*+ bl_0_205 br_0_205 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c205
*+ bl_0_205 br_0_205 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c205
*+ bl_0_205 br_0_205 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c205
*+ bl_0_205 br_0_205 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c205
*+ bl_0_205 br_0_205 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c205
*+ bl_0_205 br_0_205 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c205
*+ bl_0_205 br_0_205 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c205
*+ bl_0_205 br_0_205 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c205
*+ bl_0_205 br_0_205 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c205
*+ bl_0_205 br_0_205 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c205
*+ bl_0_205 br_0_205 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c205
*+ bl_0_205 br_0_205 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c205
*+ bl_0_205 br_0_205 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c205
*+ bl_0_205 br_0_205 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c205
*+ bl_0_205 br_0_205 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c205
*+ bl_0_205 br_0_205 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c205
*+ bl_0_205 br_0_205 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c205
*+ bl_0_205 br_0_205 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c205
*+ bl_0_205 br_0_205 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c205
*+ bl_0_205 br_0_205 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c205
*+ bl_0_205 br_0_205 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c205
*+ bl_0_205 br_0_205 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c205
*+ bl_0_205 br_0_205 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c205
*+ bl_0_205 br_0_205 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c205
*+ bl_0_205 br_0_205 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c205
*+ bl_0_205 br_0_205 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c205
*+ bl_0_205 br_0_205 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c205
*+ bl_0_205 br_0_205 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c205
*+ bl_0_205 br_0_205 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c205
*+ bl_0_205 br_0_205 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c205
*+ bl_0_205 br_0_205 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c205
*+ bl_0_205 br_0_205 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c205
*+ bl_0_205 br_0_205 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c205
*+ bl_0_205 br_0_205 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c205
*+ bl_0_205 br_0_205 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c205
*+ bl_0_205 br_0_205 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c205
*+ bl_0_205 br_0_205 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c205
*+ bl_0_205 br_0_205 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c205
*+ bl_0_205 br_0_205 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c205
*+ bl_0_205 br_0_205 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c205
*+ bl_0_205 br_0_205 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c205
*+ bl_0_205 br_0_205 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c205
*+ bl_0_205 br_0_205 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c205
*+ bl_0_205 br_0_205 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c205
*+ bl_0_205 br_0_205 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c205
*+ bl_0_205 br_0_205 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c205
*+ bl_0_205 br_0_205 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c205
*+ bl_0_205 br_0_205 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c205
*+ bl_0_205 br_0_205 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c205
*+ bl_0_205 br_0_205 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c205
*+ bl_0_205 br_0_205 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c205
*+ bl_0_205 br_0_205 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c205
*+ bl_0_205 br_0_205 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c205
*+ bl_0_205 br_0_205 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c205
*+ bl_0_205 br_0_205 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c205
*+ bl_0_205 br_0_205 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c205
*+ bl_0_205 br_0_205 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c205
*+ bl_0_205 br_0_205 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c205
*+ bl_0_205 br_0_205 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c205
*+ bl_0_205 br_0_205 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c205
*+ bl_0_205 br_0_205 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c205
*+ bl_0_205 br_0_205 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c205
*+ bl_0_205 br_0_205 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c205
*+ bl_0_205 br_0_205 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c205
*+ bl_0_205 br_0_205 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c205
*+ bl_0_205 br_0_205 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c205
*+ bl_0_205 br_0_205 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c205
*+ bl_0_205 br_0_205 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c205
*+ bl_0_205 br_0_205 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c205
*+ bl_0_205 br_0_205 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c205
*+ bl_0_205 br_0_205 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c205
*+ bl_0_205 br_0_205 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c205
*+ bl_0_205 br_0_205 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c205
*+ bl_0_205 br_0_205 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c205
*+ bl_0_205 br_0_205 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c205
*+ bl_0_205 br_0_205 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c205
*+ bl_0_205 br_0_205 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c205
*+ bl_0_205 br_0_205 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c205
*+ bl_0_205 br_0_205 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c205
*+ bl_0_205 br_0_205 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c205
*+ bl_0_205 br_0_205 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c205
*+ bl_0_205 br_0_205 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c205
*+ bl_0_205 br_0_205 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c205
*+ bl_0_205 br_0_205 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c205
*+ bl_0_205 br_0_205 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c205
*+ bl_0_205 br_0_205 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c205
*+ bl_0_205 br_0_205 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c205
*+ bl_0_205 br_0_205 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c205
*+ bl_0_205 br_0_205 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c205
*+ bl_0_205 br_0_205 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c205
*+ bl_0_205 br_0_205 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c205
*+ bl_0_205 br_0_205 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c205
*+ bl_0_205 br_0_205 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c205
*+ bl_0_205 br_0_205 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c205
*+ bl_0_205 br_0_205 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c205
*+ bl_0_205 br_0_205 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c205
*+ bl_0_205 br_0_205 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c205
*+ bl_0_205 br_0_205 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c205
*+ bl_0_205 br_0_205 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c205
*+ bl_0_205 br_0_205 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c205
*+ bl_0_205 br_0_205 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c205
*+ bl_0_205 br_0_205 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c205
*+ bl_0_205 br_0_205 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c205
*+ bl_0_205 br_0_205 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c205
*+ bl_0_205 br_0_205 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c205
*+ bl_0_205 br_0_205 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c205
*+ bl_0_205 br_0_205 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c205
*+ bl_0_205 br_0_205 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c205
*+ bl_0_205 br_0_205 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c205
+ bl_0_205 br_0_205 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c206
+ bl_0_206 br_0_206 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c206
*+ bl_0_206 br_0_206 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c206
*+ bl_0_206 br_0_206 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c206
*+ bl_0_206 br_0_206 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c206
*+ bl_0_206 br_0_206 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c206
*+ bl_0_206 br_0_206 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c206
*+ bl_0_206 br_0_206 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c206
*+ bl_0_206 br_0_206 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c206
*+ bl_0_206 br_0_206 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c206
*+ bl_0_206 br_0_206 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c206
*+ bl_0_206 br_0_206 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c206
*+ bl_0_206 br_0_206 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c206
*+ bl_0_206 br_0_206 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c206
*+ bl_0_206 br_0_206 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c206
*+ bl_0_206 br_0_206 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c206
*+ bl_0_206 br_0_206 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c206
*+ bl_0_206 br_0_206 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c206
*+ bl_0_206 br_0_206 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c206
*+ bl_0_206 br_0_206 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c206
*+ bl_0_206 br_0_206 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c206
*+ bl_0_206 br_0_206 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c206
*+ bl_0_206 br_0_206 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c206
*+ bl_0_206 br_0_206 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c206
*+ bl_0_206 br_0_206 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c206
*+ bl_0_206 br_0_206 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c206
*+ bl_0_206 br_0_206 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c206
*+ bl_0_206 br_0_206 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c206
*+ bl_0_206 br_0_206 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c206
*+ bl_0_206 br_0_206 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c206
*+ bl_0_206 br_0_206 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c206
*+ bl_0_206 br_0_206 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c206
*+ bl_0_206 br_0_206 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c206
*+ bl_0_206 br_0_206 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c206
*+ bl_0_206 br_0_206 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c206
*+ bl_0_206 br_0_206 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c206
*+ bl_0_206 br_0_206 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c206
*+ bl_0_206 br_0_206 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c206
*+ bl_0_206 br_0_206 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c206
*+ bl_0_206 br_0_206 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c206
*+ bl_0_206 br_0_206 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c206
*+ bl_0_206 br_0_206 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c206
*+ bl_0_206 br_0_206 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c206
*+ bl_0_206 br_0_206 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c206
*+ bl_0_206 br_0_206 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c206
*+ bl_0_206 br_0_206 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c206
*+ bl_0_206 br_0_206 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c206
*+ bl_0_206 br_0_206 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c206
*+ bl_0_206 br_0_206 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c206
*+ bl_0_206 br_0_206 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c206
*+ bl_0_206 br_0_206 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c206
*+ bl_0_206 br_0_206 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c206
*+ bl_0_206 br_0_206 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c206
*+ bl_0_206 br_0_206 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c206
*+ bl_0_206 br_0_206 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c206
*+ bl_0_206 br_0_206 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c206
*+ bl_0_206 br_0_206 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c206
*+ bl_0_206 br_0_206 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c206
*+ bl_0_206 br_0_206 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c206
*+ bl_0_206 br_0_206 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c206
*+ bl_0_206 br_0_206 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c206
*+ bl_0_206 br_0_206 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c206
*+ bl_0_206 br_0_206 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c206
*+ bl_0_206 br_0_206 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c206
*+ bl_0_206 br_0_206 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c206
*+ bl_0_206 br_0_206 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c206
*+ bl_0_206 br_0_206 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c206
*+ bl_0_206 br_0_206 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c206
*+ bl_0_206 br_0_206 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c206
*+ bl_0_206 br_0_206 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c206
*+ bl_0_206 br_0_206 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c206
*+ bl_0_206 br_0_206 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c206
*+ bl_0_206 br_0_206 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c206
*+ bl_0_206 br_0_206 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c206
*+ bl_0_206 br_0_206 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c206
*+ bl_0_206 br_0_206 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c206
*+ bl_0_206 br_0_206 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c206
*+ bl_0_206 br_0_206 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c206
*+ bl_0_206 br_0_206 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c206
*+ bl_0_206 br_0_206 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c206
*+ bl_0_206 br_0_206 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c206
*+ bl_0_206 br_0_206 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c206
*+ bl_0_206 br_0_206 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c206
*+ bl_0_206 br_0_206 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c206
*+ bl_0_206 br_0_206 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c206
*+ bl_0_206 br_0_206 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c206
*+ bl_0_206 br_0_206 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c206
*+ bl_0_206 br_0_206 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c206
*+ bl_0_206 br_0_206 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c206
*+ bl_0_206 br_0_206 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c206
*+ bl_0_206 br_0_206 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c206
*+ bl_0_206 br_0_206 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c206
*+ bl_0_206 br_0_206 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c206
*+ bl_0_206 br_0_206 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c206
*+ bl_0_206 br_0_206 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c206
*+ bl_0_206 br_0_206 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c206
*+ bl_0_206 br_0_206 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c206
*+ bl_0_206 br_0_206 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c206
*+ bl_0_206 br_0_206 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c206
*+ bl_0_206 br_0_206 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c206
*+ bl_0_206 br_0_206 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c206
*+ bl_0_206 br_0_206 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c206
*+ bl_0_206 br_0_206 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c206
*+ bl_0_206 br_0_206 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c206
*+ bl_0_206 br_0_206 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c206
*+ bl_0_206 br_0_206 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c206
*+ bl_0_206 br_0_206 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c206
*+ bl_0_206 br_0_206 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c206
*+ bl_0_206 br_0_206 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c206
*+ bl_0_206 br_0_206 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c206
*+ bl_0_206 br_0_206 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c206
*+ bl_0_206 br_0_206 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c206
*+ bl_0_206 br_0_206 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c206
*+ bl_0_206 br_0_206 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c206
*+ bl_0_206 br_0_206 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c206
*+ bl_0_206 br_0_206 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c206
*+ bl_0_206 br_0_206 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c206
*+ bl_0_206 br_0_206 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c206
*+ bl_0_206 br_0_206 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c206
*+ bl_0_206 br_0_206 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c206
*+ bl_0_206 br_0_206 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c206
*+ bl_0_206 br_0_206 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c206
*+ bl_0_206 br_0_206 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c206
*+ bl_0_206 br_0_206 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c206
*+ bl_0_206 br_0_206 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c206
*+ bl_0_206 br_0_206 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c206
*+ bl_0_206 br_0_206 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c206
*+ bl_0_206 br_0_206 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c206
+ bl_0_206 br_0_206 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c207
+ bl_0_207 br_0_207 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c207
*+ bl_0_207 br_0_207 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c207
*+ bl_0_207 br_0_207 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c207
*+ bl_0_207 br_0_207 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c207
*+ bl_0_207 br_0_207 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c207
*+ bl_0_207 br_0_207 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c207
*+ bl_0_207 br_0_207 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c207
*+ bl_0_207 br_0_207 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c207
*+ bl_0_207 br_0_207 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c207
*+ bl_0_207 br_0_207 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c207
*+ bl_0_207 br_0_207 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c207
*+ bl_0_207 br_0_207 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c207
*+ bl_0_207 br_0_207 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c207
*+ bl_0_207 br_0_207 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c207
*+ bl_0_207 br_0_207 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c207
*+ bl_0_207 br_0_207 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c207
*+ bl_0_207 br_0_207 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c207
*+ bl_0_207 br_0_207 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c207
*+ bl_0_207 br_0_207 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c207
*+ bl_0_207 br_0_207 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c207
*+ bl_0_207 br_0_207 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c207
*+ bl_0_207 br_0_207 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c207
*+ bl_0_207 br_0_207 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c207
*+ bl_0_207 br_0_207 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c207
*+ bl_0_207 br_0_207 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c207
*+ bl_0_207 br_0_207 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c207
*+ bl_0_207 br_0_207 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c207
*+ bl_0_207 br_0_207 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c207
*+ bl_0_207 br_0_207 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c207
*+ bl_0_207 br_0_207 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c207
*+ bl_0_207 br_0_207 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c207
*+ bl_0_207 br_0_207 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c207
*+ bl_0_207 br_0_207 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c207
*+ bl_0_207 br_0_207 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c207
*+ bl_0_207 br_0_207 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c207
*+ bl_0_207 br_0_207 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c207
*+ bl_0_207 br_0_207 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c207
*+ bl_0_207 br_0_207 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c207
*+ bl_0_207 br_0_207 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c207
*+ bl_0_207 br_0_207 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c207
*+ bl_0_207 br_0_207 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c207
*+ bl_0_207 br_0_207 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c207
*+ bl_0_207 br_0_207 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c207
*+ bl_0_207 br_0_207 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c207
*+ bl_0_207 br_0_207 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c207
*+ bl_0_207 br_0_207 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c207
*+ bl_0_207 br_0_207 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c207
*+ bl_0_207 br_0_207 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c207
*+ bl_0_207 br_0_207 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c207
*+ bl_0_207 br_0_207 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c207
*+ bl_0_207 br_0_207 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c207
*+ bl_0_207 br_0_207 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c207
*+ bl_0_207 br_0_207 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c207
*+ bl_0_207 br_0_207 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c207
*+ bl_0_207 br_0_207 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c207
*+ bl_0_207 br_0_207 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c207
*+ bl_0_207 br_0_207 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c207
*+ bl_0_207 br_0_207 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c207
*+ bl_0_207 br_0_207 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c207
*+ bl_0_207 br_0_207 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c207
*+ bl_0_207 br_0_207 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c207
*+ bl_0_207 br_0_207 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c207
*+ bl_0_207 br_0_207 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c207
*+ bl_0_207 br_0_207 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c207
*+ bl_0_207 br_0_207 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c207
*+ bl_0_207 br_0_207 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c207
*+ bl_0_207 br_0_207 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c207
*+ bl_0_207 br_0_207 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c207
*+ bl_0_207 br_0_207 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c207
*+ bl_0_207 br_0_207 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c207
*+ bl_0_207 br_0_207 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c207
*+ bl_0_207 br_0_207 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c207
*+ bl_0_207 br_0_207 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c207
*+ bl_0_207 br_0_207 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c207
*+ bl_0_207 br_0_207 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c207
*+ bl_0_207 br_0_207 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c207
*+ bl_0_207 br_0_207 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c207
*+ bl_0_207 br_0_207 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c207
*+ bl_0_207 br_0_207 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c207
*+ bl_0_207 br_0_207 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c207
*+ bl_0_207 br_0_207 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c207
*+ bl_0_207 br_0_207 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c207
*+ bl_0_207 br_0_207 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c207
*+ bl_0_207 br_0_207 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c207
*+ bl_0_207 br_0_207 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c207
*+ bl_0_207 br_0_207 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c207
*+ bl_0_207 br_0_207 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c207
*+ bl_0_207 br_0_207 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c207
*+ bl_0_207 br_0_207 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c207
*+ bl_0_207 br_0_207 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c207
*+ bl_0_207 br_0_207 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c207
*+ bl_0_207 br_0_207 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c207
*+ bl_0_207 br_0_207 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c207
*+ bl_0_207 br_0_207 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c207
*+ bl_0_207 br_0_207 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c207
*+ bl_0_207 br_0_207 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c207
*+ bl_0_207 br_0_207 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c207
*+ bl_0_207 br_0_207 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c207
*+ bl_0_207 br_0_207 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c207
*+ bl_0_207 br_0_207 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c207
*+ bl_0_207 br_0_207 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c207
*+ bl_0_207 br_0_207 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c207
*+ bl_0_207 br_0_207 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c207
*+ bl_0_207 br_0_207 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c207
*+ bl_0_207 br_0_207 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c207
*+ bl_0_207 br_0_207 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c207
*+ bl_0_207 br_0_207 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c207
*+ bl_0_207 br_0_207 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c207
*+ bl_0_207 br_0_207 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c207
*+ bl_0_207 br_0_207 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c207
*+ bl_0_207 br_0_207 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c207
*+ bl_0_207 br_0_207 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c207
*+ bl_0_207 br_0_207 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c207
*+ bl_0_207 br_0_207 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c207
*+ bl_0_207 br_0_207 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c207
*+ bl_0_207 br_0_207 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c207
*+ bl_0_207 br_0_207 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c207
*+ bl_0_207 br_0_207 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c207
*+ bl_0_207 br_0_207 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c207
*+ bl_0_207 br_0_207 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c207
*+ bl_0_207 br_0_207 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c207
*+ bl_0_207 br_0_207 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c207
*+ bl_0_207 br_0_207 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c207
*+ bl_0_207 br_0_207 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c207
*+ bl_0_207 br_0_207 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c207
*+ bl_0_207 br_0_207 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c207
*+ bl_0_207 br_0_207 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c207
+ bl_0_207 br_0_207 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c208
+ bl_0_208 br_0_208 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c208
*+ bl_0_208 br_0_208 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c208
*+ bl_0_208 br_0_208 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c208
*+ bl_0_208 br_0_208 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c208
*+ bl_0_208 br_0_208 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c208
*+ bl_0_208 br_0_208 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c208
*+ bl_0_208 br_0_208 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c208
*+ bl_0_208 br_0_208 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c208
*+ bl_0_208 br_0_208 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c208
*+ bl_0_208 br_0_208 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c208
*+ bl_0_208 br_0_208 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c208
*+ bl_0_208 br_0_208 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c208
*+ bl_0_208 br_0_208 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c208
*+ bl_0_208 br_0_208 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c208
*+ bl_0_208 br_0_208 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c208
*+ bl_0_208 br_0_208 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c208
*+ bl_0_208 br_0_208 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c208
*+ bl_0_208 br_0_208 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c208
*+ bl_0_208 br_0_208 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c208
*+ bl_0_208 br_0_208 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c208
*+ bl_0_208 br_0_208 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c208
*+ bl_0_208 br_0_208 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c208
*+ bl_0_208 br_0_208 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c208
*+ bl_0_208 br_0_208 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c208
*+ bl_0_208 br_0_208 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c208
*+ bl_0_208 br_0_208 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c208
*+ bl_0_208 br_0_208 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c208
*+ bl_0_208 br_0_208 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c208
*+ bl_0_208 br_0_208 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c208
*+ bl_0_208 br_0_208 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c208
*+ bl_0_208 br_0_208 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c208
*+ bl_0_208 br_0_208 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c208
*+ bl_0_208 br_0_208 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c208
*+ bl_0_208 br_0_208 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c208
*+ bl_0_208 br_0_208 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c208
*+ bl_0_208 br_0_208 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c208
*+ bl_0_208 br_0_208 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c208
*+ bl_0_208 br_0_208 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c208
*+ bl_0_208 br_0_208 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c208
*+ bl_0_208 br_0_208 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c208
*+ bl_0_208 br_0_208 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c208
*+ bl_0_208 br_0_208 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c208
*+ bl_0_208 br_0_208 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c208
*+ bl_0_208 br_0_208 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c208
*+ bl_0_208 br_0_208 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c208
*+ bl_0_208 br_0_208 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c208
*+ bl_0_208 br_0_208 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c208
*+ bl_0_208 br_0_208 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c208
*+ bl_0_208 br_0_208 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c208
*+ bl_0_208 br_0_208 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c208
*+ bl_0_208 br_0_208 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c208
*+ bl_0_208 br_0_208 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c208
*+ bl_0_208 br_0_208 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c208
*+ bl_0_208 br_0_208 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c208
*+ bl_0_208 br_0_208 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c208
*+ bl_0_208 br_0_208 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c208
*+ bl_0_208 br_0_208 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c208
*+ bl_0_208 br_0_208 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c208
*+ bl_0_208 br_0_208 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c208
*+ bl_0_208 br_0_208 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c208
*+ bl_0_208 br_0_208 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c208
*+ bl_0_208 br_0_208 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c208
*+ bl_0_208 br_0_208 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c208
*+ bl_0_208 br_0_208 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c208
*+ bl_0_208 br_0_208 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c208
*+ bl_0_208 br_0_208 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c208
*+ bl_0_208 br_0_208 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c208
*+ bl_0_208 br_0_208 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c208
*+ bl_0_208 br_0_208 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c208
*+ bl_0_208 br_0_208 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c208
*+ bl_0_208 br_0_208 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c208
*+ bl_0_208 br_0_208 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c208
*+ bl_0_208 br_0_208 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c208
*+ bl_0_208 br_0_208 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c208
*+ bl_0_208 br_0_208 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c208
*+ bl_0_208 br_0_208 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c208
*+ bl_0_208 br_0_208 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c208
*+ bl_0_208 br_0_208 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c208
*+ bl_0_208 br_0_208 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c208
*+ bl_0_208 br_0_208 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c208
*+ bl_0_208 br_0_208 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c208
*+ bl_0_208 br_0_208 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c208
*+ bl_0_208 br_0_208 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c208
*+ bl_0_208 br_0_208 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c208
*+ bl_0_208 br_0_208 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c208
*+ bl_0_208 br_0_208 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c208
*+ bl_0_208 br_0_208 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c208
*+ bl_0_208 br_0_208 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c208
*+ bl_0_208 br_0_208 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c208
*+ bl_0_208 br_0_208 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c208
*+ bl_0_208 br_0_208 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c208
*+ bl_0_208 br_0_208 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c208
*+ bl_0_208 br_0_208 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c208
*+ bl_0_208 br_0_208 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c208
*+ bl_0_208 br_0_208 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c208
*+ bl_0_208 br_0_208 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c208
*+ bl_0_208 br_0_208 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c208
*+ bl_0_208 br_0_208 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c208
*+ bl_0_208 br_0_208 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c208
*+ bl_0_208 br_0_208 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c208
*+ bl_0_208 br_0_208 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c208
*+ bl_0_208 br_0_208 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c208
*+ bl_0_208 br_0_208 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c208
*+ bl_0_208 br_0_208 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c208
*+ bl_0_208 br_0_208 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c208
*+ bl_0_208 br_0_208 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c208
*+ bl_0_208 br_0_208 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c208
*+ bl_0_208 br_0_208 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c208
*+ bl_0_208 br_0_208 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c208
*+ bl_0_208 br_0_208 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c208
*+ bl_0_208 br_0_208 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c208
*+ bl_0_208 br_0_208 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c208
*+ bl_0_208 br_0_208 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c208
*+ bl_0_208 br_0_208 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c208
*+ bl_0_208 br_0_208 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c208
*+ bl_0_208 br_0_208 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c208
*+ bl_0_208 br_0_208 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c208
*+ bl_0_208 br_0_208 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c208
*+ bl_0_208 br_0_208 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c208
*+ bl_0_208 br_0_208 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c208
*+ bl_0_208 br_0_208 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c208
*+ bl_0_208 br_0_208 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c208
*+ bl_0_208 br_0_208 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c208
*+ bl_0_208 br_0_208 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c208
*+ bl_0_208 br_0_208 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c208
*+ bl_0_208 br_0_208 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c208
*+ bl_0_208 br_0_208 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c208
+ bl_0_208 br_0_208 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c209
+ bl_0_209 br_0_209 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c209
*+ bl_0_209 br_0_209 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c209
*+ bl_0_209 br_0_209 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c209
*+ bl_0_209 br_0_209 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c209
*+ bl_0_209 br_0_209 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c209
*+ bl_0_209 br_0_209 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c209
*+ bl_0_209 br_0_209 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c209
*+ bl_0_209 br_0_209 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c209
*+ bl_0_209 br_0_209 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c209
*+ bl_0_209 br_0_209 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c209
*+ bl_0_209 br_0_209 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c209
*+ bl_0_209 br_0_209 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c209
*+ bl_0_209 br_0_209 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c209
*+ bl_0_209 br_0_209 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c209
*+ bl_0_209 br_0_209 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c209
*+ bl_0_209 br_0_209 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c209
*+ bl_0_209 br_0_209 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c209
*+ bl_0_209 br_0_209 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c209
*+ bl_0_209 br_0_209 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c209
*+ bl_0_209 br_0_209 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c209
*+ bl_0_209 br_0_209 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c209
*+ bl_0_209 br_0_209 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c209
*+ bl_0_209 br_0_209 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c209
*+ bl_0_209 br_0_209 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c209
*+ bl_0_209 br_0_209 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c209
*+ bl_0_209 br_0_209 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c209
*+ bl_0_209 br_0_209 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c209
*+ bl_0_209 br_0_209 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c209
*+ bl_0_209 br_0_209 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c209
*+ bl_0_209 br_0_209 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c209
*+ bl_0_209 br_0_209 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c209
*+ bl_0_209 br_0_209 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c209
*+ bl_0_209 br_0_209 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c209
*+ bl_0_209 br_0_209 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c209
*+ bl_0_209 br_0_209 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c209
*+ bl_0_209 br_0_209 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c209
*+ bl_0_209 br_0_209 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c209
*+ bl_0_209 br_0_209 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c209
*+ bl_0_209 br_0_209 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c209
*+ bl_0_209 br_0_209 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c209
*+ bl_0_209 br_0_209 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c209
*+ bl_0_209 br_0_209 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c209
*+ bl_0_209 br_0_209 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c209
*+ bl_0_209 br_0_209 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c209
*+ bl_0_209 br_0_209 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c209
*+ bl_0_209 br_0_209 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c209
*+ bl_0_209 br_0_209 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c209
*+ bl_0_209 br_0_209 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c209
*+ bl_0_209 br_0_209 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c209
*+ bl_0_209 br_0_209 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c209
*+ bl_0_209 br_0_209 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c209
*+ bl_0_209 br_0_209 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c209
*+ bl_0_209 br_0_209 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c209
*+ bl_0_209 br_0_209 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c209
*+ bl_0_209 br_0_209 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c209
*+ bl_0_209 br_0_209 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c209
*+ bl_0_209 br_0_209 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c209
*+ bl_0_209 br_0_209 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c209
*+ bl_0_209 br_0_209 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c209
*+ bl_0_209 br_0_209 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c209
*+ bl_0_209 br_0_209 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c209
*+ bl_0_209 br_0_209 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c209
*+ bl_0_209 br_0_209 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c209
*+ bl_0_209 br_0_209 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c209
*+ bl_0_209 br_0_209 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c209
*+ bl_0_209 br_0_209 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c209
*+ bl_0_209 br_0_209 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c209
*+ bl_0_209 br_0_209 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c209
*+ bl_0_209 br_0_209 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c209
*+ bl_0_209 br_0_209 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c209
*+ bl_0_209 br_0_209 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c209
*+ bl_0_209 br_0_209 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c209
*+ bl_0_209 br_0_209 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c209
*+ bl_0_209 br_0_209 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c209
*+ bl_0_209 br_0_209 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c209
*+ bl_0_209 br_0_209 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c209
*+ bl_0_209 br_0_209 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c209
*+ bl_0_209 br_0_209 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c209
*+ bl_0_209 br_0_209 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c209
*+ bl_0_209 br_0_209 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c209
*+ bl_0_209 br_0_209 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c209
*+ bl_0_209 br_0_209 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c209
*+ bl_0_209 br_0_209 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c209
*+ bl_0_209 br_0_209 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c209
*+ bl_0_209 br_0_209 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c209
*+ bl_0_209 br_0_209 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c209
*+ bl_0_209 br_0_209 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c209
*+ bl_0_209 br_0_209 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c209
*+ bl_0_209 br_0_209 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c209
*+ bl_0_209 br_0_209 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c209
*+ bl_0_209 br_0_209 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c209
*+ bl_0_209 br_0_209 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c209
*+ bl_0_209 br_0_209 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c209
*+ bl_0_209 br_0_209 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c209
*+ bl_0_209 br_0_209 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c209
*+ bl_0_209 br_0_209 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c209
*+ bl_0_209 br_0_209 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c209
*+ bl_0_209 br_0_209 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c209
*+ bl_0_209 br_0_209 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c209
*+ bl_0_209 br_0_209 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c209
*+ bl_0_209 br_0_209 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c209
*+ bl_0_209 br_0_209 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c209
*+ bl_0_209 br_0_209 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c209
*+ bl_0_209 br_0_209 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c209
*+ bl_0_209 br_0_209 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c209
*+ bl_0_209 br_0_209 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c209
*+ bl_0_209 br_0_209 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c209
*+ bl_0_209 br_0_209 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c209
*+ bl_0_209 br_0_209 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c209
*+ bl_0_209 br_0_209 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c209
*+ bl_0_209 br_0_209 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c209
*+ bl_0_209 br_0_209 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c209
*+ bl_0_209 br_0_209 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c209
*+ bl_0_209 br_0_209 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c209
*+ bl_0_209 br_0_209 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c209
*+ bl_0_209 br_0_209 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c209
*+ bl_0_209 br_0_209 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c209
*+ bl_0_209 br_0_209 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c209
*+ bl_0_209 br_0_209 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c209
*+ bl_0_209 br_0_209 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c209
*+ bl_0_209 br_0_209 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c209
*+ bl_0_209 br_0_209 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c209
*+ bl_0_209 br_0_209 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c209
*+ bl_0_209 br_0_209 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c209
*+ bl_0_209 br_0_209 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c209
*+ bl_0_209 br_0_209 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c209
*+ bl_0_209 br_0_209 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c209
+ bl_0_209 br_0_209 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c210
+ bl_0_210 br_0_210 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c210
*+ bl_0_210 br_0_210 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c210
*+ bl_0_210 br_0_210 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c210
*+ bl_0_210 br_0_210 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c210
*+ bl_0_210 br_0_210 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c210
*+ bl_0_210 br_0_210 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c210
*+ bl_0_210 br_0_210 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c210
*+ bl_0_210 br_0_210 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c210
*+ bl_0_210 br_0_210 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c210
*+ bl_0_210 br_0_210 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c210
*+ bl_0_210 br_0_210 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c210
*+ bl_0_210 br_0_210 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c210
*+ bl_0_210 br_0_210 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c210
*+ bl_0_210 br_0_210 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c210
*+ bl_0_210 br_0_210 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c210
*+ bl_0_210 br_0_210 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c210
*+ bl_0_210 br_0_210 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c210
*+ bl_0_210 br_0_210 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c210
*+ bl_0_210 br_0_210 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c210
*+ bl_0_210 br_0_210 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c210
*+ bl_0_210 br_0_210 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c210
*+ bl_0_210 br_0_210 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c210
*+ bl_0_210 br_0_210 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c210
*+ bl_0_210 br_0_210 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c210
*+ bl_0_210 br_0_210 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c210
*+ bl_0_210 br_0_210 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c210
*+ bl_0_210 br_0_210 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c210
*+ bl_0_210 br_0_210 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c210
*+ bl_0_210 br_0_210 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c210
*+ bl_0_210 br_0_210 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c210
*+ bl_0_210 br_0_210 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c210
*+ bl_0_210 br_0_210 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c210
*+ bl_0_210 br_0_210 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c210
*+ bl_0_210 br_0_210 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c210
*+ bl_0_210 br_0_210 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c210
*+ bl_0_210 br_0_210 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c210
*+ bl_0_210 br_0_210 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c210
*+ bl_0_210 br_0_210 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c210
*+ bl_0_210 br_0_210 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c210
*+ bl_0_210 br_0_210 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c210
*+ bl_0_210 br_0_210 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c210
*+ bl_0_210 br_0_210 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c210
*+ bl_0_210 br_0_210 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c210
*+ bl_0_210 br_0_210 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c210
*+ bl_0_210 br_0_210 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c210
*+ bl_0_210 br_0_210 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c210
*+ bl_0_210 br_0_210 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c210
*+ bl_0_210 br_0_210 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c210
*+ bl_0_210 br_0_210 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c210
*+ bl_0_210 br_0_210 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c210
*+ bl_0_210 br_0_210 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c210
*+ bl_0_210 br_0_210 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c210
*+ bl_0_210 br_0_210 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c210
*+ bl_0_210 br_0_210 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c210
*+ bl_0_210 br_0_210 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c210
*+ bl_0_210 br_0_210 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c210
*+ bl_0_210 br_0_210 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c210
*+ bl_0_210 br_0_210 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c210
*+ bl_0_210 br_0_210 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c210
*+ bl_0_210 br_0_210 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c210
*+ bl_0_210 br_0_210 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c210
*+ bl_0_210 br_0_210 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c210
*+ bl_0_210 br_0_210 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c210
*+ bl_0_210 br_0_210 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c210
*+ bl_0_210 br_0_210 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c210
*+ bl_0_210 br_0_210 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c210
*+ bl_0_210 br_0_210 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c210
*+ bl_0_210 br_0_210 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c210
*+ bl_0_210 br_0_210 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c210
*+ bl_0_210 br_0_210 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c210
*+ bl_0_210 br_0_210 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c210
*+ bl_0_210 br_0_210 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c210
*+ bl_0_210 br_0_210 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c210
*+ bl_0_210 br_0_210 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c210
*+ bl_0_210 br_0_210 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c210
*+ bl_0_210 br_0_210 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c210
*+ bl_0_210 br_0_210 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c210
*+ bl_0_210 br_0_210 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c210
*+ bl_0_210 br_0_210 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c210
*+ bl_0_210 br_0_210 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c210
*+ bl_0_210 br_0_210 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c210
*+ bl_0_210 br_0_210 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c210
*+ bl_0_210 br_0_210 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c210
*+ bl_0_210 br_0_210 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c210
*+ bl_0_210 br_0_210 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c210
*+ bl_0_210 br_0_210 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c210
*+ bl_0_210 br_0_210 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c210
*+ bl_0_210 br_0_210 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c210
*+ bl_0_210 br_0_210 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c210
*+ bl_0_210 br_0_210 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c210
*+ bl_0_210 br_0_210 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c210
*+ bl_0_210 br_0_210 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c210
*+ bl_0_210 br_0_210 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c210
*+ bl_0_210 br_0_210 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c210
*+ bl_0_210 br_0_210 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c210
*+ bl_0_210 br_0_210 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c210
*+ bl_0_210 br_0_210 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c210
*+ bl_0_210 br_0_210 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c210
*+ bl_0_210 br_0_210 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c210
*+ bl_0_210 br_0_210 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c210
*+ bl_0_210 br_0_210 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c210
*+ bl_0_210 br_0_210 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c210
*+ bl_0_210 br_0_210 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c210
*+ bl_0_210 br_0_210 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c210
*+ bl_0_210 br_0_210 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c210
*+ bl_0_210 br_0_210 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c210
*+ bl_0_210 br_0_210 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c210
*+ bl_0_210 br_0_210 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c210
*+ bl_0_210 br_0_210 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c210
*+ bl_0_210 br_0_210 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c210
*+ bl_0_210 br_0_210 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c210
*+ bl_0_210 br_0_210 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c210
*+ bl_0_210 br_0_210 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c210
*+ bl_0_210 br_0_210 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c210
*+ bl_0_210 br_0_210 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c210
*+ bl_0_210 br_0_210 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c210
*+ bl_0_210 br_0_210 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c210
*+ bl_0_210 br_0_210 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c210
*+ bl_0_210 br_0_210 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c210
*+ bl_0_210 br_0_210 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c210
*+ bl_0_210 br_0_210 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c210
*+ bl_0_210 br_0_210 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c210
*+ bl_0_210 br_0_210 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c210
*+ bl_0_210 br_0_210 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c210
*+ bl_0_210 br_0_210 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c210
*+ bl_0_210 br_0_210 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c210
*+ bl_0_210 br_0_210 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c210
+ bl_0_210 br_0_210 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c211
+ bl_0_211 br_0_211 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c211
*+ bl_0_211 br_0_211 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c211
*+ bl_0_211 br_0_211 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c211
*+ bl_0_211 br_0_211 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c211
*+ bl_0_211 br_0_211 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c211
*+ bl_0_211 br_0_211 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c211
*+ bl_0_211 br_0_211 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c211
*+ bl_0_211 br_0_211 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c211
*+ bl_0_211 br_0_211 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c211
*+ bl_0_211 br_0_211 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c211
*+ bl_0_211 br_0_211 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c211
*+ bl_0_211 br_0_211 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c211
*+ bl_0_211 br_0_211 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c211
*+ bl_0_211 br_0_211 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c211
*+ bl_0_211 br_0_211 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c211
*+ bl_0_211 br_0_211 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c211
*+ bl_0_211 br_0_211 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c211
*+ bl_0_211 br_0_211 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c211
*+ bl_0_211 br_0_211 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c211
*+ bl_0_211 br_0_211 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c211
*+ bl_0_211 br_0_211 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c211
*+ bl_0_211 br_0_211 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c211
*+ bl_0_211 br_0_211 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c211
*+ bl_0_211 br_0_211 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c211
*+ bl_0_211 br_0_211 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c211
*+ bl_0_211 br_0_211 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c211
*+ bl_0_211 br_0_211 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c211
*+ bl_0_211 br_0_211 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c211
*+ bl_0_211 br_0_211 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c211
*+ bl_0_211 br_0_211 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c211
*+ bl_0_211 br_0_211 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c211
*+ bl_0_211 br_0_211 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c211
*+ bl_0_211 br_0_211 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c211
*+ bl_0_211 br_0_211 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c211
*+ bl_0_211 br_0_211 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c211
*+ bl_0_211 br_0_211 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c211
*+ bl_0_211 br_0_211 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c211
*+ bl_0_211 br_0_211 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c211
*+ bl_0_211 br_0_211 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c211
*+ bl_0_211 br_0_211 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c211
*+ bl_0_211 br_0_211 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c211
*+ bl_0_211 br_0_211 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c211
*+ bl_0_211 br_0_211 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c211
*+ bl_0_211 br_0_211 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c211
*+ bl_0_211 br_0_211 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c211
*+ bl_0_211 br_0_211 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c211
*+ bl_0_211 br_0_211 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c211
*+ bl_0_211 br_0_211 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c211
*+ bl_0_211 br_0_211 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c211
*+ bl_0_211 br_0_211 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c211
*+ bl_0_211 br_0_211 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c211
*+ bl_0_211 br_0_211 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c211
*+ bl_0_211 br_0_211 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c211
*+ bl_0_211 br_0_211 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c211
*+ bl_0_211 br_0_211 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c211
*+ bl_0_211 br_0_211 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c211
*+ bl_0_211 br_0_211 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c211
*+ bl_0_211 br_0_211 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c211
*+ bl_0_211 br_0_211 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c211
*+ bl_0_211 br_0_211 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c211
*+ bl_0_211 br_0_211 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c211
*+ bl_0_211 br_0_211 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c211
*+ bl_0_211 br_0_211 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c211
*+ bl_0_211 br_0_211 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c211
*+ bl_0_211 br_0_211 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c211
*+ bl_0_211 br_0_211 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c211
*+ bl_0_211 br_0_211 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c211
*+ bl_0_211 br_0_211 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c211
*+ bl_0_211 br_0_211 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c211
*+ bl_0_211 br_0_211 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c211
*+ bl_0_211 br_0_211 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c211
*+ bl_0_211 br_0_211 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c211
*+ bl_0_211 br_0_211 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c211
*+ bl_0_211 br_0_211 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c211
*+ bl_0_211 br_0_211 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c211
*+ bl_0_211 br_0_211 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c211
*+ bl_0_211 br_0_211 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c211
*+ bl_0_211 br_0_211 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c211
*+ bl_0_211 br_0_211 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c211
*+ bl_0_211 br_0_211 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c211
*+ bl_0_211 br_0_211 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c211
*+ bl_0_211 br_0_211 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c211
*+ bl_0_211 br_0_211 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c211
*+ bl_0_211 br_0_211 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c211
*+ bl_0_211 br_0_211 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c211
*+ bl_0_211 br_0_211 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c211
*+ bl_0_211 br_0_211 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c211
*+ bl_0_211 br_0_211 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c211
*+ bl_0_211 br_0_211 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c211
*+ bl_0_211 br_0_211 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c211
*+ bl_0_211 br_0_211 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c211
*+ bl_0_211 br_0_211 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c211
*+ bl_0_211 br_0_211 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c211
*+ bl_0_211 br_0_211 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c211
*+ bl_0_211 br_0_211 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c211
*+ bl_0_211 br_0_211 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c211
*+ bl_0_211 br_0_211 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c211
*+ bl_0_211 br_0_211 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c211
*+ bl_0_211 br_0_211 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c211
*+ bl_0_211 br_0_211 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c211
*+ bl_0_211 br_0_211 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c211
*+ bl_0_211 br_0_211 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c211
*+ bl_0_211 br_0_211 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c211
*+ bl_0_211 br_0_211 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c211
*+ bl_0_211 br_0_211 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c211
*+ bl_0_211 br_0_211 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c211
*+ bl_0_211 br_0_211 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c211
*+ bl_0_211 br_0_211 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c211
*+ bl_0_211 br_0_211 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c211
*+ bl_0_211 br_0_211 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c211
*+ bl_0_211 br_0_211 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c211
*+ bl_0_211 br_0_211 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c211
*+ bl_0_211 br_0_211 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c211
*+ bl_0_211 br_0_211 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c211
*+ bl_0_211 br_0_211 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c211
*+ bl_0_211 br_0_211 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c211
*+ bl_0_211 br_0_211 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c211
*+ bl_0_211 br_0_211 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c211
*+ bl_0_211 br_0_211 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c211
*+ bl_0_211 br_0_211 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c211
*+ bl_0_211 br_0_211 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c211
*+ bl_0_211 br_0_211 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c211
*+ bl_0_211 br_0_211 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c211
*+ bl_0_211 br_0_211 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c211
*+ bl_0_211 br_0_211 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c211
*+ bl_0_211 br_0_211 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c211
*+ bl_0_211 br_0_211 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c211
+ bl_0_211 br_0_211 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c212
+ bl_0_212 br_0_212 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c212
*+ bl_0_212 br_0_212 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c212
*+ bl_0_212 br_0_212 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c212
*+ bl_0_212 br_0_212 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c212
*+ bl_0_212 br_0_212 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c212
*+ bl_0_212 br_0_212 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c212
*+ bl_0_212 br_0_212 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c212
*+ bl_0_212 br_0_212 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c212
*+ bl_0_212 br_0_212 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c212
*+ bl_0_212 br_0_212 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c212
*+ bl_0_212 br_0_212 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c212
*+ bl_0_212 br_0_212 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c212
*+ bl_0_212 br_0_212 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c212
*+ bl_0_212 br_0_212 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c212
*+ bl_0_212 br_0_212 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c212
*+ bl_0_212 br_0_212 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c212
*+ bl_0_212 br_0_212 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c212
*+ bl_0_212 br_0_212 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c212
*+ bl_0_212 br_0_212 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c212
*+ bl_0_212 br_0_212 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c212
*+ bl_0_212 br_0_212 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c212
*+ bl_0_212 br_0_212 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c212
*+ bl_0_212 br_0_212 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c212
*+ bl_0_212 br_0_212 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c212
*+ bl_0_212 br_0_212 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c212
*+ bl_0_212 br_0_212 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c212
*+ bl_0_212 br_0_212 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c212
*+ bl_0_212 br_0_212 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c212
*+ bl_0_212 br_0_212 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c212
*+ bl_0_212 br_0_212 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c212
*+ bl_0_212 br_0_212 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c212
*+ bl_0_212 br_0_212 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c212
*+ bl_0_212 br_0_212 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c212
*+ bl_0_212 br_0_212 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c212
*+ bl_0_212 br_0_212 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c212
*+ bl_0_212 br_0_212 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c212
*+ bl_0_212 br_0_212 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c212
*+ bl_0_212 br_0_212 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c212
*+ bl_0_212 br_0_212 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c212
*+ bl_0_212 br_0_212 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c212
*+ bl_0_212 br_0_212 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c212
*+ bl_0_212 br_0_212 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c212
*+ bl_0_212 br_0_212 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c212
*+ bl_0_212 br_0_212 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c212
*+ bl_0_212 br_0_212 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c212
*+ bl_0_212 br_0_212 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c212
*+ bl_0_212 br_0_212 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c212
*+ bl_0_212 br_0_212 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c212
*+ bl_0_212 br_0_212 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c212
*+ bl_0_212 br_0_212 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c212
*+ bl_0_212 br_0_212 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c212
*+ bl_0_212 br_0_212 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c212
*+ bl_0_212 br_0_212 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c212
*+ bl_0_212 br_0_212 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c212
*+ bl_0_212 br_0_212 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c212
*+ bl_0_212 br_0_212 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c212
*+ bl_0_212 br_0_212 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c212
*+ bl_0_212 br_0_212 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c212
*+ bl_0_212 br_0_212 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c212
*+ bl_0_212 br_0_212 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c212
*+ bl_0_212 br_0_212 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c212
*+ bl_0_212 br_0_212 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c212
*+ bl_0_212 br_0_212 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c212
*+ bl_0_212 br_0_212 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c212
*+ bl_0_212 br_0_212 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c212
*+ bl_0_212 br_0_212 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c212
*+ bl_0_212 br_0_212 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c212
*+ bl_0_212 br_0_212 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c212
*+ bl_0_212 br_0_212 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c212
*+ bl_0_212 br_0_212 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c212
*+ bl_0_212 br_0_212 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c212
*+ bl_0_212 br_0_212 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c212
*+ bl_0_212 br_0_212 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c212
*+ bl_0_212 br_0_212 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c212
*+ bl_0_212 br_0_212 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c212
*+ bl_0_212 br_0_212 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c212
*+ bl_0_212 br_0_212 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c212
*+ bl_0_212 br_0_212 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c212
*+ bl_0_212 br_0_212 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c212
*+ bl_0_212 br_0_212 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c212
*+ bl_0_212 br_0_212 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c212
*+ bl_0_212 br_0_212 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c212
*+ bl_0_212 br_0_212 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c212
*+ bl_0_212 br_0_212 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c212
*+ bl_0_212 br_0_212 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c212
*+ bl_0_212 br_0_212 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c212
*+ bl_0_212 br_0_212 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c212
*+ bl_0_212 br_0_212 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c212
*+ bl_0_212 br_0_212 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c212
*+ bl_0_212 br_0_212 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c212
*+ bl_0_212 br_0_212 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c212
*+ bl_0_212 br_0_212 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c212
*+ bl_0_212 br_0_212 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c212
*+ bl_0_212 br_0_212 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c212
*+ bl_0_212 br_0_212 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c212
*+ bl_0_212 br_0_212 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c212
*+ bl_0_212 br_0_212 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c212
*+ bl_0_212 br_0_212 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c212
*+ bl_0_212 br_0_212 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c212
*+ bl_0_212 br_0_212 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c212
*+ bl_0_212 br_0_212 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c212
*+ bl_0_212 br_0_212 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c212
*+ bl_0_212 br_0_212 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c212
*+ bl_0_212 br_0_212 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c212
*+ bl_0_212 br_0_212 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c212
*+ bl_0_212 br_0_212 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c212
*+ bl_0_212 br_0_212 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c212
*+ bl_0_212 br_0_212 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c212
*+ bl_0_212 br_0_212 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c212
*+ bl_0_212 br_0_212 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c212
*+ bl_0_212 br_0_212 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c212
*+ bl_0_212 br_0_212 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c212
*+ bl_0_212 br_0_212 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c212
*+ bl_0_212 br_0_212 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c212
*+ bl_0_212 br_0_212 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c212
*+ bl_0_212 br_0_212 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c212
*+ bl_0_212 br_0_212 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c212
*+ bl_0_212 br_0_212 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c212
*+ bl_0_212 br_0_212 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c212
*+ bl_0_212 br_0_212 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c212
*+ bl_0_212 br_0_212 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c212
*+ bl_0_212 br_0_212 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c212
*+ bl_0_212 br_0_212 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c212
*+ bl_0_212 br_0_212 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c212
*+ bl_0_212 br_0_212 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c212
*+ bl_0_212 br_0_212 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c212
*+ bl_0_212 br_0_212 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c212
+ bl_0_212 br_0_212 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c213
+ bl_0_213 br_0_213 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c213
*+ bl_0_213 br_0_213 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c213
*+ bl_0_213 br_0_213 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c213
*+ bl_0_213 br_0_213 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c213
*+ bl_0_213 br_0_213 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c213
*+ bl_0_213 br_0_213 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c213
*+ bl_0_213 br_0_213 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c213
*+ bl_0_213 br_0_213 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c213
*+ bl_0_213 br_0_213 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c213
*+ bl_0_213 br_0_213 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c213
*+ bl_0_213 br_0_213 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c213
*+ bl_0_213 br_0_213 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c213
*+ bl_0_213 br_0_213 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c213
*+ bl_0_213 br_0_213 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c213
*+ bl_0_213 br_0_213 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c213
*+ bl_0_213 br_0_213 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c213
*+ bl_0_213 br_0_213 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c213
*+ bl_0_213 br_0_213 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c213
*+ bl_0_213 br_0_213 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c213
*+ bl_0_213 br_0_213 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c213
*+ bl_0_213 br_0_213 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c213
*+ bl_0_213 br_0_213 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c213
*+ bl_0_213 br_0_213 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c213
*+ bl_0_213 br_0_213 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c213
*+ bl_0_213 br_0_213 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c213
*+ bl_0_213 br_0_213 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c213
*+ bl_0_213 br_0_213 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c213
*+ bl_0_213 br_0_213 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c213
*+ bl_0_213 br_0_213 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c213
*+ bl_0_213 br_0_213 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c213
*+ bl_0_213 br_0_213 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c213
*+ bl_0_213 br_0_213 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c213
*+ bl_0_213 br_0_213 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c213
*+ bl_0_213 br_0_213 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c213
*+ bl_0_213 br_0_213 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c213
*+ bl_0_213 br_0_213 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c213
*+ bl_0_213 br_0_213 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c213
*+ bl_0_213 br_0_213 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c213
*+ bl_0_213 br_0_213 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c213
*+ bl_0_213 br_0_213 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c213
*+ bl_0_213 br_0_213 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c213
*+ bl_0_213 br_0_213 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c213
*+ bl_0_213 br_0_213 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c213
*+ bl_0_213 br_0_213 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c213
*+ bl_0_213 br_0_213 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c213
*+ bl_0_213 br_0_213 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c213
*+ bl_0_213 br_0_213 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c213
*+ bl_0_213 br_0_213 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c213
*+ bl_0_213 br_0_213 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c213
*+ bl_0_213 br_0_213 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c213
*+ bl_0_213 br_0_213 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c213
*+ bl_0_213 br_0_213 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c213
*+ bl_0_213 br_0_213 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c213
*+ bl_0_213 br_0_213 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c213
*+ bl_0_213 br_0_213 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c213
*+ bl_0_213 br_0_213 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c213
*+ bl_0_213 br_0_213 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c213
*+ bl_0_213 br_0_213 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c213
*+ bl_0_213 br_0_213 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c213
*+ bl_0_213 br_0_213 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c213
*+ bl_0_213 br_0_213 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c213
*+ bl_0_213 br_0_213 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c213
*+ bl_0_213 br_0_213 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c213
*+ bl_0_213 br_0_213 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c213
*+ bl_0_213 br_0_213 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c213
*+ bl_0_213 br_0_213 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c213
*+ bl_0_213 br_0_213 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c213
*+ bl_0_213 br_0_213 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c213
*+ bl_0_213 br_0_213 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c213
*+ bl_0_213 br_0_213 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c213
*+ bl_0_213 br_0_213 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c213
*+ bl_0_213 br_0_213 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c213
*+ bl_0_213 br_0_213 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c213
*+ bl_0_213 br_0_213 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c213
*+ bl_0_213 br_0_213 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c213
*+ bl_0_213 br_0_213 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c213
*+ bl_0_213 br_0_213 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c213
*+ bl_0_213 br_0_213 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c213
*+ bl_0_213 br_0_213 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c213
*+ bl_0_213 br_0_213 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c213
*+ bl_0_213 br_0_213 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c213
*+ bl_0_213 br_0_213 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c213
*+ bl_0_213 br_0_213 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c213
*+ bl_0_213 br_0_213 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c213
*+ bl_0_213 br_0_213 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c213
*+ bl_0_213 br_0_213 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c213
*+ bl_0_213 br_0_213 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c213
*+ bl_0_213 br_0_213 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c213
*+ bl_0_213 br_0_213 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c213
*+ bl_0_213 br_0_213 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c213
*+ bl_0_213 br_0_213 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c213
*+ bl_0_213 br_0_213 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c213
*+ bl_0_213 br_0_213 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c213
*+ bl_0_213 br_0_213 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c213
*+ bl_0_213 br_0_213 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c213
*+ bl_0_213 br_0_213 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c213
*+ bl_0_213 br_0_213 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c213
*+ bl_0_213 br_0_213 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c213
*+ bl_0_213 br_0_213 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c213
*+ bl_0_213 br_0_213 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c213
*+ bl_0_213 br_0_213 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c213
*+ bl_0_213 br_0_213 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c213
*+ bl_0_213 br_0_213 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c213
*+ bl_0_213 br_0_213 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c213
*+ bl_0_213 br_0_213 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c213
*+ bl_0_213 br_0_213 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c213
*+ bl_0_213 br_0_213 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c213
*+ bl_0_213 br_0_213 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c213
*+ bl_0_213 br_0_213 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c213
*+ bl_0_213 br_0_213 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c213
*+ bl_0_213 br_0_213 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c213
*+ bl_0_213 br_0_213 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c213
*+ bl_0_213 br_0_213 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c213
*+ bl_0_213 br_0_213 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c213
*+ bl_0_213 br_0_213 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c213
*+ bl_0_213 br_0_213 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c213
*+ bl_0_213 br_0_213 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c213
*+ bl_0_213 br_0_213 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c213
*+ bl_0_213 br_0_213 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c213
*+ bl_0_213 br_0_213 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c213
*+ bl_0_213 br_0_213 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c213
*+ bl_0_213 br_0_213 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c213
*+ bl_0_213 br_0_213 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c213
*+ bl_0_213 br_0_213 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c213
*+ bl_0_213 br_0_213 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c213
*+ bl_0_213 br_0_213 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c213
*+ bl_0_213 br_0_213 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c213
+ bl_0_213 br_0_213 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c214
+ bl_0_214 br_0_214 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c214
*+ bl_0_214 br_0_214 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c214
*+ bl_0_214 br_0_214 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c214
*+ bl_0_214 br_0_214 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c214
*+ bl_0_214 br_0_214 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c214
*+ bl_0_214 br_0_214 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c214
*+ bl_0_214 br_0_214 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c214
*+ bl_0_214 br_0_214 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c214
*+ bl_0_214 br_0_214 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c214
*+ bl_0_214 br_0_214 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c214
*+ bl_0_214 br_0_214 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c214
*+ bl_0_214 br_0_214 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c214
*+ bl_0_214 br_0_214 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c214
*+ bl_0_214 br_0_214 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c214
*+ bl_0_214 br_0_214 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c214
*+ bl_0_214 br_0_214 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c214
*+ bl_0_214 br_0_214 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c214
*+ bl_0_214 br_0_214 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c214
*+ bl_0_214 br_0_214 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c214
*+ bl_0_214 br_0_214 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c214
*+ bl_0_214 br_0_214 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c214
*+ bl_0_214 br_0_214 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c214
*+ bl_0_214 br_0_214 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c214
*+ bl_0_214 br_0_214 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c214
*+ bl_0_214 br_0_214 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c214
*+ bl_0_214 br_0_214 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c214
*+ bl_0_214 br_0_214 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c214
*+ bl_0_214 br_0_214 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c214
*+ bl_0_214 br_0_214 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c214
*+ bl_0_214 br_0_214 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c214
*+ bl_0_214 br_0_214 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c214
*+ bl_0_214 br_0_214 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c214
*+ bl_0_214 br_0_214 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c214
*+ bl_0_214 br_0_214 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c214
*+ bl_0_214 br_0_214 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c214
*+ bl_0_214 br_0_214 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c214
*+ bl_0_214 br_0_214 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c214
*+ bl_0_214 br_0_214 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c214
*+ bl_0_214 br_0_214 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c214
*+ bl_0_214 br_0_214 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c214
*+ bl_0_214 br_0_214 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c214
*+ bl_0_214 br_0_214 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c214
*+ bl_0_214 br_0_214 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c214
*+ bl_0_214 br_0_214 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c214
*+ bl_0_214 br_0_214 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c214
*+ bl_0_214 br_0_214 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c214
*+ bl_0_214 br_0_214 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c214
*+ bl_0_214 br_0_214 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c214
*+ bl_0_214 br_0_214 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c214
*+ bl_0_214 br_0_214 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c214
*+ bl_0_214 br_0_214 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c214
*+ bl_0_214 br_0_214 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c214
*+ bl_0_214 br_0_214 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c214
*+ bl_0_214 br_0_214 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c214
*+ bl_0_214 br_0_214 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c214
*+ bl_0_214 br_0_214 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c214
*+ bl_0_214 br_0_214 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c214
*+ bl_0_214 br_0_214 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c214
*+ bl_0_214 br_0_214 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c214
*+ bl_0_214 br_0_214 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c214
*+ bl_0_214 br_0_214 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c214
*+ bl_0_214 br_0_214 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c214
*+ bl_0_214 br_0_214 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c214
*+ bl_0_214 br_0_214 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c214
*+ bl_0_214 br_0_214 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c214
*+ bl_0_214 br_0_214 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c214
*+ bl_0_214 br_0_214 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c214
*+ bl_0_214 br_0_214 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c214
*+ bl_0_214 br_0_214 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c214
*+ bl_0_214 br_0_214 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c214
*+ bl_0_214 br_0_214 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c214
*+ bl_0_214 br_0_214 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c214
*+ bl_0_214 br_0_214 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c214
*+ bl_0_214 br_0_214 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c214
*+ bl_0_214 br_0_214 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c214
*+ bl_0_214 br_0_214 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c214
*+ bl_0_214 br_0_214 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c214
*+ bl_0_214 br_0_214 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c214
*+ bl_0_214 br_0_214 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c214
*+ bl_0_214 br_0_214 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c214
*+ bl_0_214 br_0_214 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c214
*+ bl_0_214 br_0_214 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c214
*+ bl_0_214 br_0_214 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c214
*+ bl_0_214 br_0_214 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c214
*+ bl_0_214 br_0_214 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c214
*+ bl_0_214 br_0_214 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c214
*+ bl_0_214 br_0_214 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c214
*+ bl_0_214 br_0_214 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c214
*+ bl_0_214 br_0_214 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c214
*+ bl_0_214 br_0_214 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c214
*+ bl_0_214 br_0_214 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c214
*+ bl_0_214 br_0_214 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c214
*+ bl_0_214 br_0_214 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c214
*+ bl_0_214 br_0_214 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c214
*+ bl_0_214 br_0_214 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c214
*+ bl_0_214 br_0_214 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c214
*+ bl_0_214 br_0_214 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c214
*+ bl_0_214 br_0_214 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c214
*+ bl_0_214 br_0_214 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c214
*+ bl_0_214 br_0_214 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c214
*+ bl_0_214 br_0_214 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c214
*+ bl_0_214 br_0_214 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c214
*+ bl_0_214 br_0_214 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c214
*+ bl_0_214 br_0_214 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c214
*+ bl_0_214 br_0_214 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c214
*+ bl_0_214 br_0_214 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c214
*+ bl_0_214 br_0_214 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c214
*+ bl_0_214 br_0_214 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c214
*+ bl_0_214 br_0_214 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c214
*+ bl_0_214 br_0_214 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c214
*+ bl_0_214 br_0_214 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c214
*+ bl_0_214 br_0_214 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c214
*+ bl_0_214 br_0_214 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c214
*+ bl_0_214 br_0_214 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c214
*+ bl_0_214 br_0_214 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c214
*+ bl_0_214 br_0_214 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c214
*+ bl_0_214 br_0_214 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c214
*+ bl_0_214 br_0_214 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c214
*+ bl_0_214 br_0_214 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c214
*+ bl_0_214 br_0_214 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c214
*+ bl_0_214 br_0_214 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c214
*+ bl_0_214 br_0_214 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c214
*+ bl_0_214 br_0_214 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c214
*+ bl_0_214 br_0_214 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c214
*+ bl_0_214 br_0_214 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c214
*+ bl_0_214 br_0_214 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c214
*+ bl_0_214 br_0_214 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c214
+ bl_0_214 br_0_214 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c215
+ bl_0_215 br_0_215 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c215
*+ bl_0_215 br_0_215 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c215
*+ bl_0_215 br_0_215 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c215
*+ bl_0_215 br_0_215 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c215
*+ bl_0_215 br_0_215 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c215
*+ bl_0_215 br_0_215 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c215
*+ bl_0_215 br_0_215 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c215
*+ bl_0_215 br_0_215 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c215
*+ bl_0_215 br_0_215 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c215
*+ bl_0_215 br_0_215 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c215
*+ bl_0_215 br_0_215 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c215
*+ bl_0_215 br_0_215 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c215
*+ bl_0_215 br_0_215 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c215
*+ bl_0_215 br_0_215 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c215
*+ bl_0_215 br_0_215 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c215
*+ bl_0_215 br_0_215 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c215
*+ bl_0_215 br_0_215 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c215
*+ bl_0_215 br_0_215 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c215
*+ bl_0_215 br_0_215 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c215
*+ bl_0_215 br_0_215 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c215
*+ bl_0_215 br_0_215 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c215
*+ bl_0_215 br_0_215 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c215
*+ bl_0_215 br_0_215 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c215
*+ bl_0_215 br_0_215 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c215
*+ bl_0_215 br_0_215 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c215
*+ bl_0_215 br_0_215 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c215
*+ bl_0_215 br_0_215 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c215
*+ bl_0_215 br_0_215 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c215
*+ bl_0_215 br_0_215 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c215
*+ bl_0_215 br_0_215 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c215
*+ bl_0_215 br_0_215 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c215
*+ bl_0_215 br_0_215 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c215
*+ bl_0_215 br_0_215 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c215
*+ bl_0_215 br_0_215 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c215
*+ bl_0_215 br_0_215 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c215
*+ bl_0_215 br_0_215 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c215
*+ bl_0_215 br_0_215 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c215
*+ bl_0_215 br_0_215 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c215
*+ bl_0_215 br_0_215 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c215
*+ bl_0_215 br_0_215 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c215
*+ bl_0_215 br_0_215 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c215
*+ bl_0_215 br_0_215 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c215
*+ bl_0_215 br_0_215 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c215
*+ bl_0_215 br_0_215 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c215
*+ bl_0_215 br_0_215 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c215
*+ bl_0_215 br_0_215 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c215
*+ bl_0_215 br_0_215 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c215
*+ bl_0_215 br_0_215 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c215
*+ bl_0_215 br_0_215 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c215
*+ bl_0_215 br_0_215 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c215
*+ bl_0_215 br_0_215 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c215
*+ bl_0_215 br_0_215 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c215
*+ bl_0_215 br_0_215 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c215
*+ bl_0_215 br_0_215 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c215
*+ bl_0_215 br_0_215 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c215
*+ bl_0_215 br_0_215 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c215
*+ bl_0_215 br_0_215 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c215
*+ bl_0_215 br_0_215 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c215
*+ bl_0_215 br_0_215 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c215
*+ bl_0_215 br_0_215 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c215
*+ bl_0_215 br_0_215 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c215
*+ bl_0_215 br_0_215 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c215
*+ bl_0_215 br_0_215 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c215
*+ bl_0_215 br_0_215 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c215
*+ bl_0_215 br_0_215 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c215
*+ bl_0_215 br_0_215 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c215
*+ bl_0_215 br_0_215 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c215
*+ bl_0_215 br_0_215 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c215
*+ bl_0_215 br_0_215 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c215
*+ bl_0_215 br_0_215 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c215
*+ bl_0_215 br_0_215 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c215
*+ bl_0_215 br_0_215 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c215
*+ bl_0_215 br_0_215 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c215
*+ bl_0_215 br_0_215 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c215
*+ bl_0_215 br_0_215 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c215
*+ bl_0_215 br_0_215 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c215
*+ bl_0_215 br_0_215 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c215
*+ bl_0_215 br_0_215 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c215
*+ bl_0_215 br_0_215 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c215
*+ bl_0_215 br_0_215 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c215
*+ bl_0_215 br_0_215 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c215
*+ bl_0_215 br_0_215 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c215
*+ bl_0_215 br_0_215 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c215
*+ bl_0_215 br_0_215 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c215
*+ bl_0_215 br_0_215 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c215
*+ bl_0_215 br_0_215 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c215
*+ bl_0_215 br_0_215 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c215
*+ bl_0_215 br_0_215 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c215
*+ bl_0_215 br_0_215 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c215
*+ bl_0_215 br_0_215 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c215
*+ bl_0_215 br_0_215 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c215
*+ bl_0_215 br_0_215 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c215
*+ bl_0_215 br_0_215 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c215
*+ bl_0_215 br_0_215 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c215
*+ bl_0_215 br_0_215 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c215
*+ bl_0_215 br_0_215 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c215
*+ bl_0_215 br_0_215 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c215
*+ bl_0_215 br_0_215 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c215
*+ bl_0_215 br_0_215 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c215
*+ bl_0_215 br_0_215 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c215
*+ bl_0_215 br_0_215 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c215
*+ bl_0_215 br_0_215 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c215
*+ bl_0_215 br_0_215 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c215
*+ bl_0_215 br_0_215 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c215
*+ bl_0_215 br_0_215 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c215
*+ bl_0_215 br_0_215 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c215
*+ bl_0_215 br_0_215 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c215
*+ bl_0_215 br_0_215 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c215
*+ bl_0_215 br_0_215 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c215
*+ bl_0_215 br_0_215 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c215
*+ bl_0_215 br_0_215 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c215
*+ bl_0_215 br_0_215 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c215
*+ bl_0_215 br_0_215 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c215
*+ bl_0_215 br_0_215 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c215
*+ bl_0_215 br_0_215 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c215
*+ bl_0_215 br_0_215 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c215
*+ bl_0_215 br_0_215 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c215
*+ bl_0_215 br_0_215 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c215
*+ bl_0_215 br_0_215 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c215
*+ bl_0_215 br_0_215 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c215
*+ bl_0_215 br_0_215 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c215
*+ bl_0_215 br_0_215 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c215
*+ bl_0_215 br_0_215 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c215
*+ bl_0_215 br_0_215 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c215
*+ bl_0_215 br_0_215 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c215
*+ bl_0_215 br_0_215 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c215
*+ bl_0_215 br_0_215 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c215
+ bl_0_215 br_0_215 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c216
+ bl_0_216 br_0_216 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c216
*+ bl_0_216 br_0_216 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c216
*+ bl_0_216 br_0_216 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c216
*+ bl_0_216 br_0_216 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c216
*+ bl_0_216 br_0_216 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c216
*+ bl_0_216 br_0_216 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c216
*+ bl_0_216 br_0_216 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c216
*+ bl_0_216 br_0_216 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c216
*+ bl_0_216 br_0_216 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c216
*+ bl_0_216 br_0_216 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c216
*+ bl_0_216 br_0_216 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c216
*+ bl_0_216 br_0_216 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c216
*+ bl_0_216 br_0_216 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c216
*+ bl_0_216 br_0_216 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c216
*+ bl_0_216 br_0_216 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c216
*+ bl_0_216 br_0_216 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c216
*+ bl_0_216 br_0_216 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c216
*+ bl_0_216 br_0_216 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c216
*+ bl_0_216 br_0_216 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c216
*+ bl_0_216 br_0_216 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c216
*+ bl_0_216 br_0_216 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c216
*+ bl_0_216 br_0_216 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c216
*+ bl_0_216 br_0_216 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c216
*+ bl_0_216 br_0_216 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c216
*+ bl_0_216 br_0_216 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c216
*+ bl_0_216 br_0_216 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c216
*+ bl_0_216 br_0_216 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c216
*+ bl_0_216 br_0_216 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c216
*+ bl_0_216 br_0_216 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c216
*+ bl_0_216 br_0_216 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c216
*+ bl_0_216 br_0_216 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c216
*+ bl_0_216 br_0_216 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c216
*+ bl_0_216 br_0_216 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c216
*+ bl_0_216 br_0_216 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c216
*+ bl_0_216 br_0_216 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c216
*+ bl_0_216 br_0_216 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c216
*+ bl_0_216 br_0_216 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c216
*+ bl_0_216 br_0_216 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c216
*+ bl_0_216 br_0_216 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c216
*+ bl_0_216 br_0_216 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c216
*+ bl_0_216 br_0_216 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c216
*+ bl_0_216 br_0_216 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c216
*+ bl_0_216 br_0_216 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c216
*+ bl_0_216 br_0_216 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c216
*+ bl_0_216 br_0_216 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c216
*+ bl_0_216 br_0_216 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c216
*+ bl_0_216 br_0_216 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c216
*+ bl_0_216 br_0_216 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c216
*+ bl_0_216 br_0_216 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c216
*+ bl_0_216 br_0_216 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c216
*+ bl_0_216 br_0_216 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c216
*+ bl_0_216 br_0_216 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c216
*+ bl_0_216 br_0_216 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c216
*+ bl_0_216 br_0_216 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c216
*+ bl_0_216 br_0_216 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c216
*+ bl_0_216 br_0_216 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c216
*+ bl_0_216 br_0_216 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c216
*+ bl_0_216 br_0_216 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c216
*+ bl_0_216 br_0_216 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c216
*+ bl_0_216 br_0_216 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c216
*+ bl_0_216 br_0_216 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c216
*+ bl_0_216 br_0_216 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c216
*+ bl_0_216 br_0_216 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c216
*+ bl_0_216 br_0_216 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c216
*+ bl_0_216 br_0_216 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c216
*+ bl_0_216 br_0_216 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c216
*+ bl_0_216 br_0_216 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c216
*+ bl_0_216 br_0_216 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c216
*+ bl_0_216 br_0_216 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c216
*+ bl_0_216 br_0_216 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c216
*+ bl_0_216 br_0_216 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c216
*+ bl_0_216 br_0_216 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c216
*+ bl_0_216 br_0_216 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c216
*+ bl_0_216 br_0_216 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c216
*+ bl_0_216 br_0_216 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c216
*+ bl_0_216 br_0_216 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c216
*+ bl_0_216 br_0_216 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c216
*+ bl_0_216 br_0_216 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c216
*+ bl_0_216 br_0_216 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c216
*+ bl_0_216 br_0_216 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c216
*+ bl_0_216 br_0_216 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c216
*+ bl_0_216 br_0_216 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c216
*+ bl_0_216 br_0_216 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c216
*+ bl_0_216 br_0_216 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c216
*+ bl_0_216 br_0_216 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c216
*+ bl_0_216 br_0_216 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c216
*+ bl_0_216 br_0_216 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c216
*+ bl_0_216 br_0_216 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c216
*+ bl_0_216 br_0_216 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c216
*+ bl_0_216 br_0_216 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c216
*+ bl_0_216 br_0_216 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c216
*+ bl_0_216 br_0_216 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c216
*+ bl_0_216 br_0_216 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c216
*+ bl_0_216 br_0_216 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c216
*+ bl_0_216 br_0_216 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c216
*+ bl_0_216 br_0_216 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c216
*+ bl_0_216 br_0_216 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c216
*+ bl_0_216 br_0_216 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c216
*+ bl_0_216 br_0_216 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c216
*+ bl_0_216 br_0_216 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c216
*+ bl_0_216 br_0_216 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c216
*+ bl_0_216 br_0_216 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c216
*+ bl_0_216 br_0_216 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c216
*+ bl_0_216 br_0_216 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c216
*+ bl_0_216 br_0_216 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c216
*+ bl_0_216 br_0_216 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c216
*+ bl_0_216 br_0_216 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c216
*+ bl_0_216 br_0_216 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c216
*+ bl_0_216 br_0_216 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c216
*+ bl_0_216 br_0_216 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c216
*+ bl_0_216 br_0_216 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c216
*+ bl_0_216 br_0_216 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c216
*+ bl_0_216 br_0_216 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c216
*+ bl_0_216 br_0_216 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c216
*+ bl_0_216 br_0_216 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c216
*+ bl_0_216 br_0_216 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c216
*+ bl_0_216 br_0_216 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c216
*+ bl_0_216 br_0_216 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c216
*+ bl_0_216 br_0_216 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c216
*+ bl_0_216 br_0_216 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c216
*+ bl_0_216 br_0_216 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c216
*+ bl_0_216 br_0_216 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c216
*+ bl_0_216 br_0_216 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c216
*+ bl_0_216 br_0_216 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c216
*+ bl_0_216 br_0_216 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c216
*+ bl_0_216 br_0_216 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c216
*+ bl_0_216 br_0_216 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c216
+ bl_0_216 br_0_216 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c217
+ bl_0_217 br_0_217 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c217
*+ bl_0_217 br_0_217 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c217
*+ bl_0_217 br_0_217 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c217
*+ bl_0_217 br_0_217 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c217
*+ bl_0_217 br_0_217 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c217
*+ bl_0_217 br_0_217 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c217
*+ bl_0_217 br_0_217 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c217
*+ bl_0_217 br_0_217 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c217
*+ bl_0_217 br_0_217 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c217
*+ bl_0_217 br_0_217 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c217
*+ bl_0_217 br_0_217 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c217
*+ bl_0_217 br_0_217 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c217
*+ bl_0_217 br_0_217 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c217
*+ bl_0_217 br_0_217 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c217
*+ bl_0_217 br_0_217 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c217
*+ bl_0_217 br_0_217 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c217
*+ bl_0_217 br_0_217 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c217
*+ bl_0_217 br_0_217 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c217
*+ bl_0_217 br_0_217 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c217
*+ bl_0_217 br_0_217 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c217
*+ bl_0_217 br_0_217 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c217
*+ bl_0_217 br_0_217 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c217
*+ bl_0_217 br_0_217 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c217
*+ bl_0_217 br_0_217 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c217
*+ bl_0_217 br_0_217 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c217
*+ bl_0_217 br_0_217 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c217
*+ bl_0_217 br_0_217 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c217
*+ bl_0_217 br_0_217 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c217
*+ bl_0_217 br_0_217 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c217
*+ bl_0_217 br_0_217 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c217
*+ bl_0_217 br_0_217 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c217
*+ bl_0_217 br_0_217 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c217
*+ bl_0_217 br_0_217 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c217
*+ bl_0_217 br_0_217 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c217
*+ bl_0_217 br_0_217 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c217
*+ bl_0_217 br_0_217 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c217
*+ bl_0_217 br_0_217 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c217
*+ bl_0_217 br_0_217 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c217
*+ bl_0_217 br_0_217 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c217
*+ bl_0_217 br_0_217 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c217
*+ bl_0_217 br_0_217 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c217
*+ bl_0_217 br_0_217 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c217
*+ bl_0_217 br_0_217 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c217
*+ bl_0_217 br_0_217 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c217
*+ bl_0_217 br_0_217 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c217
*+ bl_0_217 br_0_217 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c217
*+ bl_0_217 br_0_217 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c217
*+ bl_0_217 br_0_217 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c217
*+ bl_0_217 br_0_217 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c217
*+ bl_0_217 br_0_217 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c217
*+ bl_0_217 br_0_217 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c217
*+ bl_0_217 br_0_217 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c217
*+ bl_0_217 br_0_217 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c217
*+ bl_0_217 br_0_217 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c217
*+ bl_0_217 br_0_217 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c217
*+ bl_0_217 br_0_217 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c217
*+ bl_0_217 br_0_217 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c217
*+ bl_0_217 br_0_217 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c217
*+ bl_0_217 br_0_217 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c217
*+ bl_0_217 br_0_217 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c217
*+ bl_0_217 br_0_217 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c217
*+ bl_0_217 br_0_217 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c217
*+ bl_0_217 br_0_217 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c217
*+ bl_0_217 br_0_217 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c217
*+ bl_0_217 br_0_217 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c217
*+ bl_0_217 br_0_217 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c217
*+ bl_0_217 br_0_217 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c217
*+ bl_0_217 br_0_217 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c217
*+ bl_0_217 br_0_217 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c217
*+ bl_0_217 br_0_217 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c217
*+ bl_0_217 br_0_217 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c217
*+ bl_0_217 br_0_217 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c217
*+ bl_0_217 br_0_217 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c217
*+ bl_0_217 br_0_217 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c217
*+ bl_0_217 br_0_217 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c217
*+ bl_0_217 br_0_217 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c217
*+ bl_0_217 br_0_217 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c217
*+ bl_0_217 br_0_217 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c217
*+ bl_0_217 br_0_217 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c217
*+ bl_0_217 br_0_217 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c217
*+ bl_0_217 br_0_217 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c217
*+ bl_0_217 br_0_217 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c217
*+ bl_0_217 br_0_217 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c217
*+ bl_0_217 br_0_217 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c217
*+ bl_0_217 br_0_217 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c217
*+ bl_0_217 br_0_217 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c217
*+ bl_0_217 br_0_217 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c217
*+ bl_0_217 br_0_217 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c217
*+ bl_0_217 br_0_217 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c217
*+ bl_0_217 br_0_217 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c217
*+ bl_0_217 br_0_217 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c217
*+ bl_0_217 br_0_217 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c217
*+ bl_0_217 br_0_217 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c217
*+ bl_0_217 br_0_217 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c217
*+ bl_0_217 br_0_217 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c217
*+ bl_0_217 br_0_217 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c217
*+ bl_0_217 br_0_217 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c217
*+ bl_0_217 br_0_217 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c217
*+ bl_0_217 br_0_217 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c217
*+ bl_0_217 br_0_217 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c217
*+ bl_0_217 br_0_217 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c217
*+ bl_0_217 br_0_217 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c217
*+ bl_0_217 br_0_217 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c217
*+ bl_0_217 br_0_217 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c217
*+ bl_0_217 br_0_217 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c217
*+ bl_0_217 br_0_217 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c217
*+ bl_0_217 br_0_217 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c217
*+ bl_0_217 br_0_217 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c217
*+ bl_0_217 br_0_217 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c217
*+ bl_0_217 br_0_217 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c217
*+ bl_0_217 br_0_217 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c217
*+ bl_0_217 br_0_217 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c217
*+ bl_0_217 br_0_217 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c217
*+ bl_0_217 br_0_217 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c217
*+ bl_0_217 br_0_217 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c217
*+ bl_0_217 br_0_217 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c217
*+ bl_0_217 br_0_217 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c217
*+ bl_0_217 br_0_217 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c217
*+ bl_0_217 br_0_217 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c217
*+ bl_0_217 br_0_217 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c217
*+ bl_0_217 br_0_217 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c217
*+ bl_0_217 br_0_217 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c217
*+ bl_0_217 br_0_217 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c217
*+ bl_0_217 br_0_217 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c217
*+ bl_0_217 br_0_217 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c217
*+ bl_0_217 br_0_217 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c217
*+ bl_0_217 br_0_217 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c217
+ bl_0_217 br_0_217 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c218
+ bl_0_218 br_0_218 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c218
*+ bl_0_218 br_0_218 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c218
*+ bl_0_218 br_0_218 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c218
*+ bl_0_218 br_0_218 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c218
*+ bl_0_218 br_0_218 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c218
*+ bl_0_218 br_0_218 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c218
*+ bl_0_218 br_0_218 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c218
*+ bl_0_218 br_0_218 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c218
*+ bl_0_218 br_0_218 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c218
*+ bl_0_218 br_0_218 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c218
*+ bl_0_218 br_0_218 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c218
*+ bl_0_218 br_0_218 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c218
*+ bl_0_218 br_0_218 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c218
*+ bl_0_218 br_0_218 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c218
*+ bl_0_218 br_0_218 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c218
*+ bl_0_218 br_0_218 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c218
*+ bl_0_218 br_0_218 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c218
*+ bl_0_218 br_0_218 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c218
*+ bl_0_218 br_0_218 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c218
*+ bl_0_218 br_0_218 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c218
*+ bl_0_218 br_0_218 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c218
*+ bl_0_218 br_0_218 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c218
*+ bl_0_218 br_0_218 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c218
*+ bl_0_218 br_0_218 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c218
*+ bl_0_218 br_0_218 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c218
*+ bl_0_218 br_0_218 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c218
*+ bl_0_218 br_0_218 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c218
*+ bl_0_218 br_0_218 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c218
*+ bl_0_218 br_0_218 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c218
*+ bl_0_218 br_0_218 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c218
*+ bl_0_218 br_0_218 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c218
*+ bl_0_218 br_0_218 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c218
*+ bl_0_218 br_0_218 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c218
*+ bl_0_218 br_0_218 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c218
*+ bl_0_218 br_0_218 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c218
*+ bl_0_218 br_0_218 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c218
*+ bl_0_218 br_0_218 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c218
*+ bl_0_218 br_0_218 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c218
*+ bl_0_218 br_0_218 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c218
*+ bl_0_218 br_0_218 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c218
*+ bl_0_218 br_0_218 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c218
*+ bl_0_218 br_0_218 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c218
*+ bl_0_218 br_0_218 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c218
*+ bl_0_218 br_0_218 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c218
*+ bl_0_218 br_0_218 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c218
*+ bl_0_218 br_0_218 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c218
*+ bl_0_218 br_0_218 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c218
*+ bl_0_218 br_0_218 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c218
*+ bl_0_218 br_0_218 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c218
*+ bl_0_218 br_0_218 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c218
*+ bl_0_218 br_0_218 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c218
*+ bl_0_218 br_0_218 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c218
*+ bl_0_218 br_0_218 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c218
*+ bl_0_218 br_0_218 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c218
*+ bl_0_218 br_0_218 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c218
*+ bl_0_218 br_0_218 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c218
*+ bl_0_218 br_0_218 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c218
*+ bl_0_218 br_0_218 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c218
*+ bl_0_218 br_0_218 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c218
*+ bl_0_218 br_0_218 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c218
*+ bl_0_218 br_0_218 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c218
*+ bl_0_218 br_0_218 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c218
*+ bl_0_218 br_0_218 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c218
*+ bl_0_218 br_0_218 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c218
*+ bl_0_218 br_0_218 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c218
*+ bl_0_218 br_0_218 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c218
*+ bl_0_218 br_0_218 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c218
*+ bl_0_218 br_0_218 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c218
*+ bl_0_218 br_0_218 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c218
*+ bl_0_218 br_0_218 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c218
*+ bl_0_218 br_0_218 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c218
*+ bl_0_218 br_0_218 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c218
*+ bl_0_218 br_0_218 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c218
*+ bl_0_218 br_0_218 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c218
*+ bl_0_218 br_0_218 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c218
*+ bl_0_218 br_0_218 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c218
*+ bl_0_218 br_0_218 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c218
*+ bl_0_218 br_0_218 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c218
*+ bl_0_218 br_0_218 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c218
*+ bl_0_218 br_0_218 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c218
*+ bl_0_218 br_0_218 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c218
*+ bl_0_218 br_0_218 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c218
*+ bl_0_218 br_0_218 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c218
*+ bl_0_218 br_0_218 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c218
*+ bl_0_218 br_0_218 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c218
*+ bl_0_218 br_0_218 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c218
*+ bl_0_218 br_0_218 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c218
*+ bl_0_218 br_0_218 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c218
*+ bl_0_218 br_0_218 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c218
*+ bl_0_218 br_0_218 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c218
*+ bl_0_218 br_0_218 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c218
*+ bl_0_218 br_0_218 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c218
*+ bl_0_218 br_0_218 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c218
*+ bl_0_218 br_0_218 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c218
*+ bl_0_218 br_0_218 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c218
*+ bl_0_218 br_0_218 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c218
*+ bl_0_218 br_0_218 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c218
*+ bl_0_218 br_0_218 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c218
*+ bl_0_218 br_0_218 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c218
*+ bl_0_218 br_0_218 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c218
*+ bl_0_218 br_0_218 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c218
*+ bl_0_218 br_0_218 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c218
*+ bl_0_218 br_0_218 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c218
*+ bl_0_218 br_0_218 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c218
*+ bl_0_218 br_0_218 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c218
*+ bl_0_218 br_0_218 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c218
*+ bl_0_218 br_0_218 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c218
*+ bl_0_218 br_0_218 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c218
*+ bl_0_218 br_0_218 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c218
*+ bl_0_218 br_0_218 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c218
*+ bl_0_218 br_0_218 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c218
*+ bl_0_218 br_0_218 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c218
*+ bl_0_218 br_0_218 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c218
*+ bl_0_218 br_0_218 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c218
*+ bl_0_218 br_0_218 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c218
*+ bl_0_218 br_0_218 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c218
*+ bl_0_218 br_0_218 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c218
*+ bl_0_218 br_0_218 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c218
*+ bl_0_218 br_0_218 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c218
*+ bl_0_218 br_0_218 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c218
*+ bl_0_218 br_0_218 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c218
*+ bl_0_218 br_0_218 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c218
*+ bl_0_218 br_0_218 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c218
*+ bl_0_218 br_0_218 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c218
*+ bl_0_218 br_0_218 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c218
*+ bl_0_218 br_0_218 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c218
*+ bl_0_218 br_0_218 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c218
+ bl_0_218 br_0_218 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c219
+ bl_0_219 br_0_219 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c219
*+ bl_0_219 br_0_219 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c219
*+ bl_0_219 br_0_219 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c219
*+ bl_0_219 br_0_219 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c219
*+ bl_0_219 br_0_219 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c219
*+ bl_0_219 br_0_219 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c219
*+ bl_0_219 br_0_219 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c219
*+ bl_0_219 br_0_219 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c219
*+ bl_0_219 br_0_219 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c219
*+ bl_0_219 br_0_219 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c219
*+ bl_0_219 br_0_219 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c219
*+ bl_0_219 br_0_219 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c219
*+ bl_0_219 br_0_219 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c219
*+ bl_0_219 br_0_219 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c219
*+ bl_0_219 br_0_219 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c219
*+ bl_0_219 br_0_219 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c219
*+ bl_0_219 br_0_219 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c219
*+ bl_0_219 br_0_219 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c219
*+ bl_0_219 br_0_219 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c219
*+ bl_0_219 br_0_219 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c219
*+ bl_0_219 br_0_219 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c219
*+ bl_0_219 br_0_219 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c219
*+ bl_0_219 br_0_219 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c219
*+ bl_0_219 br_0_219 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c219
*+ bl_0_219 br_0_219 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c219
*+ bl_0_219 br_0_219 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c219
*+ bl_0_219 br_0_219 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c219
*+ bl_0_219 br_0_219 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c219
*+ bl_0_219 br_0_219 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c219
*+ bl_0_219 br_0_219 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c219
*+ bl_0_219 br_0_219 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c219
*+ bl_0_219 br_0_219 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c219
*+ bl_0_219 br_0_219 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c219
*+ bl_0_219 br_0_219 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c219
*+ bl_0_219 br_0_219 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c219
*+ bl_0_219 br_0_219 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c219
*+ bl_0_219 br_0_219 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c219
*+ bl_0_219 br_0_219 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c219
*+ bl_0_219 br_0_219 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c219
*+ bl_0_219 br_0_219 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c219
*+ bl_0_219 br_0_219 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c219
*+ bl_0_219 br_0_219 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c219
*+ bl_0_219 br_0_219 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c219
*+ bl_0_219 br_0_219 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c219
*+ bl_0_219 br_0_219 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c219
*+ bl_0_219 br_0_219 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c219
*+ bl_0_219 br_0_219 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c219
*+ bl_0_219 br_0_219 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c219
*+ bl_0_219 br_0_219 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c219
*+ bl_0_219 br_0_219 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c219
*+ bl_0_219 br_0_219 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c219
*+ bl_0_219 br_0_219 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c219
*+ bl_0_219 br_0_219 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c219
*+ bl_0_219 br_0_219 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c219
*+ bl_0_219 br_0_219 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c219
*+ bl_0_219 br_0_219 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c219
*+ bl_0_219 br_0_219 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c219
*+ bl_0_219 br_0_219 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c219
*+ bl_0_219 br_0_219 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c219
*+ bl_0_219 br_0_219 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c219
*+ bl_0_219 br_0_219 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c219
*+ bl_0_219 br_0_219 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c219
*+ bl_0_219 br_0_219 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c219
*+ bl_0_219 br_0_219 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c219
*+ bl_0_219 br_0_219 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c219
*+ bl_0_219 br_0_219 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c219
*+ bl_0_219 br_0_219 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c219
*+ bl_0_219 br_0_219 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c219
*+ bl_0_219 br_0_219 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c219
*+ bl_0_219 br_0_219 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c219
*+ bl_0_219 br_0_219 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c219
*+ bl_0_219 br_0_219 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c219
*+ bl_0_219 br_0_219 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c219
*+ bl_0_219 br_0_219 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c219
*+ bl_0_219 br_0_219 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c219
*+ bl_0_219 br_0_219 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c219
*+ bl_0_219 br_0_219 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c219
*+ bl_0_219 br_0_219 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c219
*+ bl_0_219 br_0_219 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c219
*+ bl_0_219 br_0_219 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c219
*+ bl_0_219 br_0_219 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c219
*+ bl_0_219 br_0_219 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c219
*+ bl_0_219 br_0_219 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c219
*+ bl_0_219 br_0_219 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c219
*+ bl_0_219 br_0_219 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c219
*+ bl_0_219 br_0_219 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c219
*+ bl_0_219 br_0_219 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c219
*+ bl_0_219 br_0_219 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c219
*+ bl_0_219 br_0_219 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c219
*+ bl_0_219 br_0_219 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c219
*+ bl_0_219 br_0_219 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c219
*+ bl_0_219 br_0_219 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c219
*+ bl_0_219 br_0_219 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c219
*+ bl_0_219 br_0_219 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c219
*+ bl_0_219 br_0_219 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c219
*+ bl_0_219 br_0_219 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c219
*+ bl_0_219 br_0_219 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c219
*+ bl_0_219 br_0_219 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c219
*+ bl_0_219 br_0_219 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c219
*+ bl_0_219 br_0_219 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c219
*+ bl_0_219 br_0_219 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c219
*+ bl_0_219 br_0_219 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c219
*+ bl_0_219 br_0_219 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c219
*+ bl_0_219 br_0_219 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c219
*+ bl_0_219 br_0_219 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c219
*+ bl_0_219 br_0_219 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c219
*+ bl_0_219 br_0_219 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c219
*+ bl_0_219 br_0_219 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c219
*+ bl_0_219 br_0_219 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c219
*+ bl_0_219 br_0_219 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c219
*+ bl_0_219 br_0_219 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c219
*+ bl_0_219 br_0_219 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c219
*+ bl_0_219 br_0_219 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c219
*+ bl_0_219 br_0_219 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c219
*+ bl_0_219 br_0_219 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c219
*+ bl_0_219 br_0_219 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c219
*+ bl_0_219 br_0_219 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c219
*+ bl_0_219 br_0_219 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c219
*+ bl_0_219 br_0_219 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c219
*+ bl_0_219 br_0_219 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c219
*+ bl_0_219 br_0_219 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c219
*+ bl_0_219 br_0_219 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c219
*+ bl_0_219 br_0_219 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c219
*+ bl_0_219 br_0_219 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c219
*+ bl_0_219 br_0_219 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c219
*+ bl_0_219 br_0_219 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c219
*+ bl_0_219 br_0_219 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c219
+ bl_0_219 br_0_219 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c220
+ bl_0_220 br_0_220 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c220
*+ bl_0_220 br_0_220 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c220
*+ bl_0_220 br_0_220 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c220
*+ bl_0_220 br_0_220 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c220
*+ bl_0_220 br_0_220 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c220
*+ bl_0_220 br_0_220 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c220
*+ bl_0_220 br_0_220 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c220
*+ bl_0_220 br_0_220 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c220
*+ bl_0_220 br_0_220 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c220
*+ bl_0_220 br_0_220 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c220
*+ bl_0_220 br_0_220 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c220
*+ bl_0_220 br_0_220 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c220
*+ bl_0_220 br_0_220 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c220
*+ bl_0_220 br_0_220 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c220
*+ bl_0_220 br_0_220 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c220
*+ bl_0_220 br_0_220 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c220
*+ bl_0_220 br_0_220 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c220
*+ bl_0_220 br_0_220 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c220
*+ bl_0_220 br_0_220 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c220
*+ bl_0_220 br_0_220 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c220
*+ bl_0_220 br_0_220 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c220
*+ bl_0_220 br_0_220 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c220
*+ bl_0_220 br_0_220 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c220
*+ bl_0_220 br_0_220 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c220
*+ bl_0_220 br_0_220 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c220
*+ bl_0_220 br_0_220 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c220
*+ bl_0_220 br_0_220 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c220
*+ bl_0_220 br_0_220 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c220
*+ bl_0_220 br_0_220 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c220
*+ bl_0_220 br_0_220 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c220
*+ bl_0_220 br_0_220 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c220
*+ bl_0_220 br_0_220 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c220
*+ bl_0_220 br_0_220 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c220
*+ bl_0_220 br_0_220 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c220
*+ bl_0_220 br_0_220 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c220
*+ bl_0_220 br_0_220 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c220
*+ bl_0_220 br_0_220 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c220
*+ bl_0_220 br_0_220 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c220
*+ bl_0_220 br_0_220 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c220
*+ bl_0_220 br_0_220 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c220
*+ bl_0_220 br_0_220 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c220
*+ bl_0_220 br_0_220 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c220
*+ bl_0_220 br_0_220 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c220
*+ bl_0_220 br_0_220 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c220
*+ bl_0_220 br_0_220 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c220
*+ bl_0_220 br_0_220 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c220
*+ bl_0_220 br_0_220 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c220
*+ bl_0_220 br_0_220 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c220
*+ bl_0_220 br_0_220 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c220
*+ bl_0_220 br_0_220 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c220
*+ bl_0_220 br_0_220 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c220
*+ bl_0_220 br_0_220 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c220
*+ bl_0_220 br_0_220 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c220
*+ bl_0_220 br_0_220 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c220
*+ bl_0_220 br_0_220 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c220
*+ bl_0_220 br_0_220 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c220
*+ bl_0_220 br_0_220 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c220
*+ bl_0_220 br_0_220 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c220
*+ bl_0_220 br_0_220 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c220
*+ bl_0_220 br_0_220 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c220
*+ bl_0_220 br_0_220 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c220
*+ bl_0_220 br_0_220 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c220
*+ bl_0_220 br_0_220 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c220
*+ bl_0_220 br_0_220 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c220
*+ bl_0_220 br_0_220 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c220
*+ bl_0_220 br_0_220 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c220
*+ bl_0_220 br_0_220 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c220
*+ bl_0_220 br_0_220 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c220
*+ bl_0_220 br_0_220 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c220
*+ bl_0_220 br_0_220 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c220
*+ bl_0_220 br_0_220 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c220
*+ bl_0_220 br_0_220 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c220
*+ bl_0_220 br_0_220 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c220
*+ bl_0_220 br_0_220 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c220
*+ bl_0_220 br_0_220 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c220
*+ bl_0_220 br_0_220 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c220
*+ bl_0_220 br_0_220 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c220
*+ bl_0_220 br_0_220 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c220
*+ bl_0_220 br_0_220 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c220
*+ bl_0_220 br_0_220 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c220
*+ bl_0_220 br_0_220 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c220
*+ bl_0_220 br_0_220 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c220
*+ bl_0_220 br_0_220 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c220
*+ bl_0_220 br_0_220 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c220
*+ bl_0_220 br_0_220 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c220
*+ bl_0_220 br_0_220 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c220
*+ bl_0_220 br_0_220 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c220
*+ bl_0_220 br_0_220 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c220
*+ bl_0_220 br_0_220 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c220
*+ bl_0_220 br_0_220 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c220
*+ bl_0_220 br_0_220 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c220
*+ bl_0_220 br_0_220 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c220
*+ bl_0_220 br_0_220 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c220
*+ bl_0_220 br_0_220 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c220
*+ bl_0_220 br_0_220 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c220
*+ bl_0_220 br_0_220 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c220
*+ bl_0_220 br_0_220 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c220
*+ bl_0_220 br_0_220 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c220
*+ bl_0_220 br_0_220 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c220
*+ bl_0_220 br_0_220 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c220
*+ bl_0_220 br_0_220 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c220
*+ bl_0_220 br_0_220 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c220
*+ bl_0_220 br_0_220 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c220
*+ bl_0_220 br_0_220 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c220
*+ bl_0_220 br_0_220 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c220
*+ bl_0_220 br_0_220 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c220
*+ bl_0_220 br_0_220 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c220
*+ bl_0_220 br_0_220 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c220
*+ bl_0_220 br_0_220 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c220
*+ bl_0_220 br_0_220 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c220
*+ bl_0_220 br_0_220 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c220
*+ bl_0_220 br_0_220 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c220
*+ bl_0_220 br_0_220 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c220
*+ bl_0_220 br_0_220 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c220
*+ bl_0_220 br_0_220 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c220
*+ bl_0_220 br_0_220 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c220
*+ bl_0_220 br_0_220 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c220
*+ bl_0_220 br_0_220 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c220
*+ bl_0_220 br_0_220 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c220
*+ bl_0_220 br_0_220 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c220
*+ bl_0_220 br_0_220 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c220
*+ bl_0_220 br_0_220 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c220
*+ bl_0_220 br_0_220 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c220
*+ bl_0_220 br_0_220 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c220
*+ bl_0_220 br_0_220 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c220
*+ bl_0_220 br_0_220 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c220
*+ bl_0_220 br_0_220 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c220
+ bl_0_220 br_0_220 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c221
+ bl_0_221 br_0_221 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c221
*+ bl_0_221 br_0_221 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c221
*+ bl_0_221 br_0_221 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c221
*+ bl_0_221 br_0_221 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c221
*+ bl_0_221 br_0_221 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c221
*+ bl_0_221 br_0_221 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c221
*+ bl_0_221 br_0_221 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c221
*+ bl_0_221 br_0_221 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c221
*+ bl_0_221 br_0_221 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c221
*+ bl_0_221 br_0_221 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c221
*+ bl_0_221 br_0_221 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c221
*+ bl_0_221 br_0_221 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c221
*+ bl_0_221 br_0_221 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c221
*+ bl_0_221 br_0_221 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c221
*+ bl_0_221 br_0_221 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c221
*+ bl_0_221 br_0_221 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c221
*+ bl_0_221 br_0_221 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c221
*+ bl_0_221 br_0_221 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c221
*+ bl_0_221 br_0_221 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c221
*+ bl_0_221 br_0_221 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c221
*+ bl_0_221 br_0_221 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c221
*+ bl_0_221 br_0_221 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c221
*+ bl_0_221 br_0_221 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c221
*+ bl_0_221 br_0_221 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c221
*+ bl_0_221 br_0_221 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c221
*+ bl_0_221 br_0_221 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c221
*+ bl_0_221 br_0_221 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c221
*+ bl_0_221 br_0_221 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c221
*+ bl_0_221 br_0_221 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c221
*+ bl_0_221 br_0_221 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c221
*+ bl_0_221 br_0_221 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c221
*+ bl_0_221 br_0_221 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c221
*+ bl_0_221 br_0_221 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c221
*+ bl_0_221 br_0_221 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c221
*+ bl_0_221 br_0_221 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c221
*+ bl_0_221 br_0_221 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c221
*+ bl_0_221 br_0_221 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c221
*+ bl_0_221 br_0_221 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c221
*+ bl_0_221 br_0_221 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c221
*+ bl_0_221 br_0_221 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c221
*+ bl_0_221 br_0_221 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c221
*+ bl_0_221 br_0_221 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c221
*+ bl_0_221 br_0_221 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c221
*+ bl_0_221 br_0_221 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c221
*+ bl_0_221 br_0_221 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c221
*+ bl_0_221 br_0_221 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c221
*+ bl_0_221 br_0_221 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c221
*+ bl_0_221 br_0_221 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c221
*+ bl_0_221 br_0_221 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c221
*+ bl_0_221 br_0_221 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c221
*+ bl_0_221 br_0_221 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c221
*+ bl_0_221 br_0_221 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c221
*+ bl_0_221 br_0_221 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c221
*+ bl_0_221 br_0_221 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c221
*+ bl_0_221 br_0_221 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c221
*+ bl_0_221 br_0_221 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c221
*+ bl_0_221 br_0_221 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c221
*+ bl_0_221 br_0_221 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c221
*+ bl_0_221 br_0_221 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c221
*+ bl_0_221 br_0_221 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c221
*+ bl_0_221 br_0_221 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c221
*+ bl_0_221 br_0_221 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c221
*+ bl_0_221 br_0_221 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c221
*+ bl_0_221 br_0_221 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c221
*+ bl_0_221 br_0_221 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c221
*+ bl_0_221 br_0_221 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c221
*+ bl_0_221 br_0_221 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c221
*+ bl_0_221 br_0_221 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c221
*+ bl_0_221 br_0_221 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c221
*+ bl_0_221 br_0_221 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c221
*+ bl_0_221 br_0_221 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c221
*+ bl_0_221 br_0_221 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c221
*+ bl_0_221 br_0_221 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c221
*+ bl_0_221 br_0_221 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c221
*+ bl_0_221 br_0_221 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c221
*+ bl_0_221 br_0_221 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c221
*+ bl_0_221 br_0_221 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c221
*+ bl_0_221 br_0_221 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c221
*+ bl_0_221 br_0_221 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c221
*+ bl_0_221 br_0_221 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c221
*+ bl_0_221 br_0_221 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c221
*+ bl_0_221 br_0_221 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c221
*+ bl_0_221 br_0_221 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c221
*+ bl_0_221 br_0_221 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c221
*+ bl_0_221 br_0_221 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c221
*+ bl_0_221 br_0_221 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c221
*+ bl_0_221 br_0_221 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c221
*+ bl_0_221 br_0_221 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c221
*+ bl_0_221 br_0_221 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c221
*+ bl_0_221 br_0_221 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c221
*+ bl_0_221 br_0_221 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c221
*+ bl_0_221 br_0_221 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c221
*+ bl_0_221 br_0_221 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c221
*+ bl_0_221 br_0_221 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c221
*+ bl_0_221 br_0_221 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c221
*+ bl_0_221 br_0_221 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c221
*+ bl_0_221 br_0_221 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c221
*+ bl_0_221 br_0_221 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c221
*+ bl_0_221 br_0_221 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c221
*+ bl_0_221 br_0_221 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c221
*+ bl_0_221 br_0_221 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c221
*+ bl_0_221 br_0_221 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c221
*+ bl_0_221 br_0_221 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c221
*+ bl_0_221 br_0_221 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c221
*+ bl_0_221 br_0_221 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c221
*+ bl_0_221 br_0_221 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c221
*+ bl_0_221 br_0_221 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c221
*+ bl_0_221 br_0_221 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c221
*+ bl_0_221 br_0_221 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c221
*+ bl_0_221 br_0_221 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c221
*+ bl_0_221 br_0_221 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c221
*+ bl_0_221 br_0_221 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c221
*+ bl_0_221 br_0_221 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c221
*+ bl_0_221 br_0_221 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c221
*+ bl_0_221 br_0_221 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c221
*+ bl_0_221 br_0_221 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c221
*+ bl_0_221 br_0_221 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c221
*+ bl_0_221 br_0_221 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c221
*+ bl_0_221 br_0_221 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c221
*+ bl_0_221 br_0_221 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c221
*+ bl_0_221 br_0_221 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c221
*+ bl_0_221 br_0_221 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c221
*+ bl_0_221 br_0_221 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c221
*+ bl_0_221 br_0_221 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c221
*+ bl_0_221 br_0_221 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c221
*+ bl_0_221 br_0_221 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c221
*+ bl_0_221 br_0_221 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c221
+ bl_0_221 br_0_221 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c222
+ bl_0_222 br_0_222 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c222
*+ bl_0_222 br_0_222 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c222
*+ bl_0_222 br_0_222 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c222
*+ bl_0_222 br_0_222 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c222
*+ bl_0_222 br_0_222 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c222
*+ bl_0_222 br_0_222 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c222
*+ bl_0_222 br_0_222 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c222
*+ bl_0_222 br_0_222 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c222
*+ bl_0_222 br_0_222 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c222
*+ bl_0_222 br_0_222 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c222
*+ bl_0_222 br_0_222 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c222
*+ bl_0_222 br_0_222 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c222
*+ bl_0_222 br_0_222 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c222
*+ bl_0_222 br_0_222 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c222
*+ bl_0_222 br_0_222 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c222
*+ bl_0_222 br_0_222 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c222
*+ bl_0_222 br_0_222 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c222
*+ bl_0_222 br_0_222 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c222
*+ bl_0_222 br_0_222 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c222
*+ bl_0_222 br_0_222 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c222
*+ bl_0_222 br_0_222 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c222
*+ bl_0_222 br_0_222 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c222
*+ bl_0_222 br_0_222 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c222
*+ bl_0_222 br_0_222 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c222
*+ bl_0_222 br_0_222 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c222
*+ bl_0_222 br_0_222 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c222
*+ bl_0_222 br_0_222 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c222
*+ bl_0_222 br_0_222 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c222
*+ bl_0_222 br_0_222 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c222
*+ bl_0_222 br_0_222 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c222
*+ bl_0_222 br_0_222 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c222
*+ bl_0_222 br_0_222 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c222
*+ bl_0_222 br_0_222 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c222
*+ bl_0_222 br_0_222 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c222
*+ bl_0_222 br_0_222 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c222
*+ bl_0_222 br_0_222 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c222
*+ bl_0_222 br_0_222 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c222
*+ bl_0_222 br_0_222 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c222
*+ bl_0_222 br_0_222 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c222
*+ bl_0_222 br_0_222 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c222
*+ bl_0_222 br_0_222 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c222
*+ bl_0_222 br_0_222 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c222
*+ bl_0_222 br_0_222 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c222
*+ bl_0_222 br_0_222 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c222
*+ bl_0_222 br_0_222 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c222
*+ bl_0_222 br_0_222 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c222
*+ bl_0_222 br_0_222 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c222
*+ bl_0_222 br_0_222 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c222
*+ bl_0_222 br_0_222 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c222
*+ bl_0_222 br_0_222 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c222
*+ bl_0_222 br_0_222 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c222
*+ bl_0_222 br_0_222 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c222
*+ bl_0_222 br_0_222 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c222
*+ bl_0_222 br_0_222 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c222
*+ bl_0_222 br_0_222 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c222
*+ bl_0_222 br_0_222 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c222
*+ bl_0_222 br_0_222 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c222
*+ bl_0_222 br_0_222 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c222
*+ bl_0_222 br_0_222 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c222
*+ bl_0_222 br_0_222 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c222
*+ bl_0_222 br_0_222 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c222
*+ bl_0_222 br_0_222 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c222
*+ bl_0_222 br_0_222 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c222
*+ bl_0_222 br_0_222 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c222
*+ bl_0_222 br_0_222 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c222
*+ bl_0_222 br_0_222 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c222
*+ bl_0_222 br_0_222 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c222
*+ bl_0_222 br_0_222 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c222
*+ bl_0_222 br_0_222 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c222
*+ bl_0_222 br_0_222 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c222
*+ bl_0_222 br_0_222 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c222
*+ bl_0_222 br_0_222 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c222
*+ bl_0_222 br_0_222 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c222
*+ bl_0_222 br_0_222 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c222
*+ bl_0_222 br_0_222 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c222
*+ bl_0_222 br_0_222 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c222
*+ bl_0_222 br_0_222 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c222
*+ bl_0_222 br_0_222 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c222
*+ bl_0_222 br_0_222 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c222
*+ bl_0_222 br_0_222 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c222
*+ bl_0_222 br_0_222 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c222
*+ bl_0_222 br_0_222 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c222
*+ bl_0_222 br_0_222 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c222
*+ bl_0_222 br_0_222 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c222
*+ bl_0_222 br_0_222 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c222
*+ bl_0_222 br_0_222 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c222
*+ bl_0_222 br_0_222 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c222
*+ bl_0_222 br_0_222 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c222
*+ bl_0_222 br_0_222 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c222
*+ bl_0_222 br_0_222 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c222
*+ bl_0_222 br_0_222 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c222
*+ bl_0_222 br_0_222 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c222
*+ bl_0_222 br_0_222 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c222
*+ bl_0_222 br_0_222 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c222
*+ bl_0_222 br_0_222 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c222
*+ bl_0_222 br_0_222 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c222
*+ bl_0_222 br_0_222 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c222
*+ bl_0_222 br_0_222 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c222
*+ bl_0_222 br_0_222 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c222
*+ bl_0_222 br_0_222 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c222
*+ bl_0_222 br_0_222 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c222
*+ bl_0_222 br_0_222 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c222
*+ bl_0_222 br_0_222 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c222
*+ bl_0_222 br_0_222 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c222
*+ bl_0_222 br_0_222 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c222
*+ bl_0_222 br_0_222 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c222
*+ bl_0_222 br_0_222 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c222
*+ bl_0_222 br_0_222 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c222
*+ bl_0_222 br_0_222 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c222
*+ bl_0_222 br_0_222 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c222
*+ bl_0_222 br_0_222 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c222
*+ bl_0_222 br_0_222 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c222
*+ bl_0_222 br_0_222 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c222
*+ bl_0_222 br_0_222 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c222
*+ bl_0_222 br_0_222 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c222
*+ bl_0_222 br_0_222 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c222
*+ bl_0_222 br_0_222 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c222
*+ bl_0_222 br_0_222 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c222
*+ bl_0_222 br_0_222 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c222
*+ bl_0_222 br_0_222 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c222
*+ bl_0_222 br_0_222 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c222
*+ bl_0_222 br_0_222 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c222
*+ bl_0_222 br_0_222 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c222
*+ bl_0_222 br_0_222 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c222
*+ bl_0_222 br_0_222 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c222
*+ bl_0_222 br_0_222 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c222
*+ bl_0_222 br_0_222 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c222
+ bl_0_222 br_0_222 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c223
+ bl_0_223 br_0_223 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c223
*+ bl_0_223 br_0_223 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c223
*+ bl_0_223 br_0_223 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c223
*+ bl_0_223 br_0_223 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c223
*+ bl_0_223 br_0_223 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c223
*+ bl_0_223 br_0_223 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c223
*+ bl_0_223 br_0_223 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c223
*+ bl_0_223 br_0_223 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c223
*+ bl_0_223 br_0_223 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c223
*+ bl_0_223 br_0_223 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c223
*+ bl_0_223 br_0_223 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c223
*+ bl_0_223 br_0_223 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c223
*+ bl_0_223 br_0_223 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c223
*+ bl_0_223 br_0_223 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c223
*+ bl_0_223 br_0_223 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c223
*+ bl_0_223 br_0_223 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c223
*+ bl_0_223 br_0_223 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c223
*+ bl_0_223 br_0_223 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c223
*+ bl_0_223 br_0_223 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c223
*+ bl_0_223 br_0_223 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c223
*+ bl_0_223 br_0_223 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c223
*+ bl_0_223 br_0_223 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c223
*+ bl_0_223 br_0_223 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c223
*+ bl_0_223 br_0_223 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c223
*+ bl_0_223 br_0_223 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c223
*+ bl_0_223 br_0_223 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c223
*+ bl_0_223 br_0_223 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c223
*+ bl_0_223 br_0_223 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c223
*+ bl_0_223 br_0_223 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c223
*+ bl_0_223 br_0_223 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c223
*+ bl_0_223 br_0_223 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c223
*+ bl_0_223 br_0_223 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c223
*+ bl_0_223 br_0_223 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c223
*+ bl_0_223 br_0_223 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c223
*+ bl_0_223 br_0_223 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c223
*+ bl_0_223 br_0_223 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c223
*+ bl_0_223 br_0_223 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c223
*+ bl_0_223 br_0_223 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c223
*+ bl_0_223 br_0_223 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c223
*+ bl_0_223 br_0_223 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c223
*+ bl_0_223 br_0_223 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c223
*+ bl_0_223 br_0_223 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c223
*+ bl_0_223 br_0_223 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c223
*+ bl_0_223 br_0_223 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c223
*+ bl_0_223 br_0_223 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c223
*+ bl_0_223 br_0_223 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c223
*+ bl_0_223 br_0_223 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c223
*+ bl_0_223 br_0_223 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c223
*+ bl_0_223 br_0_223 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c223
*+ bl_0_223 br_0_223 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c223
*+ bl_0_223 br_0_223 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c223
*+ bl_0_223 br_0_223 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c223
*+ bl_0_223 br_0_223 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c223
*+ bl_0_223 br_0_223 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c223
*+ bl_0_223 br_0_223 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c223
*+ bl_0_223 br_0_223 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c223
*+ bl_0_223 br_0_223 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c223
*+ bl_0_223 br_0_223 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c223
*+ bl_0_223 br_0_223 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c223
*+ bl_0_223 br_0_223 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c223
*+ bl_0_223 br_0_223 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c223
*+ bl_0_223 br_0_223 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c223
*+ bl_0_223 br_0_223 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c223
*+ bl_0_223 br_0_223 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c223
*+ bl_0_223 br_0_223 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c223
*+ bl_0_223 br_0_223 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c223
*+ bl_0_223 br_0_223 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c223
*+ bl_0_223 br_0_223 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c223
*+ bl_0_223 br_0_223 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c223
*+ bl_0_223 br_0_223 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c223
*+ bl_0_223 br_0_223 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c223
*+ bl_0_223 br_0_223 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c223
*+ bl_0_223 br_0_223 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c223
*+ bl_0_223 br_0_223 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c223
*+ bl_0_223 br_0_223 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c223
*+ bl_0_223 br_0_223 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c223
*+ bl_0_223 br_0_223 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c223
*+ bl_0_223 br_0_223 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c223
*+ bl_0_223 br_0_223 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c223
*+ bl_0_223 br_0_223 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c223
*+ bl_0_223 br_0_223 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c223
*+ bl_0_223 br_0_223 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c223
*+ bl_0_223 br_0_223 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c223
*+ bl_0_223 br_0_223 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c223
*+ bl_0_223 br_0_223 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c223
*+ bl_0_223 br_0_223 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c223
*+ bl_0_223 br_0_223 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c223
*+ bl_0_223 br_0_223 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c223
*+ bl_0_223 br_0_223 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c223
*+ bl_0_223 br_0_223 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c223
*+ bl_0_223 br_0_223 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c223
*+ bl_0_223 br_0_223 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c223
*+ bl_0_223 br_0_223 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c223
*+ bl_0_223 br_0_223 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c223
*+ bl_0_223 br_0_223 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c223
*+ bl_0_223 br_0_223 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c223
*+ bl_0_223 br_0_223 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c223
*+ bl_0_223 br_0_223 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c223
*+ bl_0_223 br_0_223 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c223
*+ bl_0_223 br_0_223 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c223
*+ bl_0_223 br_0_223 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c223
*+ bl_0_223 br_0_223 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c223
*+ bl_0_223 br_0_223 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c223
*+ bl_0_223 br_0_223 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c223
*+ bl_0_223 br_0_223 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c223
*+ bl_0_223 br_0_223 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c223
*+ bl_0_223 br_0_223 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c223
*+ bl_0_223 br_0_223 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c223
*+ bl_0_223 br_0_223 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c223
*+ bl_0_223 br_0_223 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c223
*+ bl_0_223 br_0_223 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c223
*+ bl_0_223 br_0_223 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c223
*+ bl_0_223 br_0_223 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c223
*+ bl_0_223 br_0_223 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c223
*+ bl_0_223 br_0_223 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c223
*+ bl_0_223 br_0_223 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c223
*+ bl_0_223 br_0_223 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c223
*+ bl_0_223 br_0_223 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c223
*+ bl_0_223 br_0_223 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c223
*+ bl_0_223 br_0_223 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c223
*+ bl_0_223 br_0_223 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c223
*+ bl_0_223 br_0_223 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c223
*+ bl_0_223 br_0_223 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c223
*+ bl_0_223 br_0_223 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c223
*+ bl_0_223 br_0_223 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c223
*+ bl_0_223 br_0_223 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c223
*+ bl_0_223 br_0_223 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c223
+ bl_0_223 br_0_223 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c224
+ bl_0_224 br_0_224 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c224
*+ bl_0_224 br_0_224 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c224
*+ bl_0_224 br_0_224 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c224
*+ bl_0_224 br_0_224 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c224
*+ bl_0_224 br_0_224 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c224
*+ bl_0_224 br_0_224 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c224
*+ bl_0_224 br_0_224 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c224
*+ bl_0_224 br_0_224 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c224
*+ bl_0_224 br_0_224 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c224
*+ bl_0_224 br_0_224 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c224
*+ bl_0_224 br_0_224 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c224
*+ bl_0_224 br_0_224 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c224
*+ bl_0_224 br_0_224 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c224
*+ bl_0_224 br_0_224 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c224
*+ bl_0_224 br_0_224 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c224
*+ bl_0_224 br_0_224 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c224
*+ bl_0_224 br_0_224 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c224
*+ bl_0_224 br_0_224 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c224
*+ bl_0_224 br_0_224 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c224
*+ bl_0_224 br_0_224 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c224
*+ bl_0_224 br_0_224 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c224
*+ bl_0_224 br_0_224 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c224
*+ bl_0_224 br_0_224 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c224
*+ bl_0_224 br_0_224 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c224
*+ bl_0_224 br_0_224 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c224
*+ bl_0_224 br_0_224 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c224
*+ bl_0_224 br_0_224 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c224
*+ bl_0_224 br_0_224 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c224
*+ bl_0_224 br_0_224 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c224
*+ bl_0_224 br_0_224 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c224
*+ bl_0_224 br_0_224 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c224
*+ bl_0_224 br_0_224 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c224
*+ bl_0_224 br_0_224 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c224
*+ bl_0_224 br_0_224 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c224
*+ bl_0_224 br_0_224 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c224
*+ bl_0_224 br_0_224 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c224
*+ bl_0_224 br_0_224 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c224
*+ bl_0_224 br_0_224 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c224
*+ bl_0_224 br_0_224 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c224
*+ bl_0_224 br_0_224 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c224
*+ bl_0_224 br_0_224 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c224
*+ bl_0_224 br_0_224 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c224
*+ bl_0_224 br_0_224 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c224
*+ bl_0_224 br_0_224 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c224
*+ bl_0_224 br_0_224 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c224
*+ bl_0_224 br_0_224 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c224
*+ bl_0_224 br_0_224 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c224
*+ bl_0_224 br_0_224 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c224
*+ bl_0_224 br_0_224 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c224
*+ bl_0_224 br_0_224 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c224
*+ bl_0_224 br_0_224 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c224
*+ bl_0_224 br_0_224 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c224
*+ bl_0_224 br_0_224 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c224
*+ bl_0_224 br_0_224 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c224
*+ bl_0_224 br_0_224 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c224
*+ bl_0_224 br_0_224 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c224
*+ bl_0_224 br_0_224 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c224
*+ bl_0_224 br_0_224 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c224
*+ bl_0_224 br_0_224 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c224
*+ bl_0_224 br_0_224 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c224
*+ bl_0_224 br_0_224 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c224
*+ bl_0_224 br_0_224 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c224
*+ bl_0_224 br_0_224 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c224
*+ bl_0_224 br_0_224 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c224
*+ bl_0_224 br_0_224 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c224
*+ bl_0_224 br_0_224 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c224
*+ bl_0_224 br_0_224 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c224
*+ bl_0_224 br_0_224 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c224
*+ bl_0_224 br_0_224 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c224
*+ bl_0_224 br_0_224 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c224
*+ bl_0_224 br_0_224 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c224
*+ bl_0_224 br_0_224 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c224
*+ bl_0_224 br_0_224 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c224
*+ bl_0_224 br_0_224 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c224
*+ bl_0_224 br_0_224 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c224
*+ bl_0_224 br_0_224 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c224
*+ bl_0_224 br_0_224 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c224
*+ bl_0_224 br_0_224 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c224
*+ bl_0_224 br_0_224 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c224
*+ bl_0_224 br_0_224 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c224
*+ bl_0_224 br_0_224 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c224
*+ bl_0_224 br_0_224 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c224
*+ bl_0_224 br_0_224 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c224
*+ bl_0_224 br_0_224 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c224
*+ bl_0_224 br_0_224 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c224
*+ bl_0_224 br_0_224 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c224
*+ bl_0_224 br_0_224 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c224
*+ bl_0_224 br_0_224 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c224
*+ bl_0_224 br_0_224 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c224
*+ bl_0_224 br_0_224 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c224
*+ bl_0_224 br_0_224 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c224
*+ bl_0_224 br_0_224 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c224
*+ bl_0_224 br_0_224 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c224
*+ bl_0_224 br_0_224 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c224
*+ bl_0_224 br_0_224 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c224
*+ bl_0_224 br_0_224 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c224
*+ bl_0_224 br_0_224 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c224
*+ bl_0_224 br_0_224 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c224
*+ bl_0_224 br_0_224 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c224
*+ bl_0_224 br_0_224 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c224
*+ bl_0_224 br_0_224 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c224
*+ bl_0_224 br_0_224 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c224
*+ bl_0_224 br_0_224 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c224
*+ bl_0_224 br_0_224 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c224
*+ bl_0_224 br_0_224 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c224
*+ bl_0_224 br_0_224 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c224
*+ bl_0_224 br_0_224 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c224
*+ bl_0_224 br_0_224 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c224
*+ bl_0_224 br_0_224 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c224
*+ bl_0_224 br_0_224 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c224
*+ bl_0_224 br_0_224 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c224
*+ bl_0_224 br_0_224 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c224
*+ bl_0_224 br_0_224 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c224
*+ bl_0_224 br_0_224 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c224
*+ bl_0_224 br_0_224 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c224
*+ bl_0_224 br_0_224 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c224
*+ bl_0_224 br_0_224 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c224
*+ bl_0_224 br_0_224 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c224
*+ bl_0_224 br_0_224 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c224
*+ bl_0_224 br_0_224 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c224
*+ bl_0_224 br_0_224 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c224
*+ bl_0_224 br_0_224 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c224
*+ bl_0_224 br_0_224 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c224
*+ bl_0_224 br_0_224 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c224
*+ bl_0_224 br_0_224 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c224
*+ bl_0_224 br_0_224 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c224
*+ bl_0_224 br_0_224 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c224
+ bl_0_224 br_0_224 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c225
+ bl_0_225 br_0_225 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c225
*+ bl_0_225 br_0_225 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c225
*+ bl_0_225 br_0_225 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c225
*+ bl_0_225 br_0_225 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c225
*+ bl_0_225 br_0_225 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c225
*+ bl_0_225 br_0_225 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c225
*+ bl_0_225 br_0_225 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c225
*+ bl_0_225 br_0_225 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c225
*+ bl_0_225 br_0_225 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c225
*+ bl_0_225 br_0_225 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c225
*+ bl_0_225 br_0_225 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c225
*+ bl_0_225 br_0_225 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c225
*+ bl_0_225 br_0_225 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c225
*+ bl_0_225 br_0_225 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c225
*+ bl_0_225 br_0_225 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c225
*+ bl_0_225 br_0_225 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c225
*+ bl_0_225 br_0_225 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c225
*+ bl_0_225 br_0_225 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c225
*+ bl_0_225 br_0_225 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c225
*+ bl_0_225 br_0_225 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c225
*+ bl_0_225 br_0_225 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c225
*+ bl_0_225 br_0_225 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c225
*+ bl_0_225 br_0_225 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c225
*+ bl_0_225 br_0_225 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c225
*+ bl_0_225 br_0_225 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c225
*+ bl_0_225 br_0_225 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c225
*+ bl_0_225 br_0_225 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c225
*+ bl_0_225 br_0_225 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c225
*+ bl_0_225 br_0_225 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c225
*+ bl_0_225 br_0_225 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c225
*+ bl_0_225 br_0_225 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c225
*+ bl_0_225 br_0_225 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c225
*+ bl_0_225 br_0_225 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c225
*+ bl_0_225 br_0_225 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c225
*+ bl_0_225 br_0_225 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c225
*+ bl_0_225 br_0_225 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c225
*+ bl_0_225 br_0_225 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c225
*+ bl_0_225 br_0_225 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c225
*+ bl_0_225 br_0_225 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c225
*+ bl_0_225 br_0_225 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c225
*+ bl_0_225 br_0_225 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c225
*+ bl_0_225 br_0_225 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c225
*+ bl_0_225 br_0_225 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c225
*+ bl_0_225 br_0_225 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c225
*+ bl_0_225 br_0_225 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c225
*+ bl_0_225 br_0_225 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c225
*+ bl_0_225 br_0_225 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c225
*+ bl_0_225 br_0_225 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c225
*+ bl_0_225 br_0_225 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c225
*+ bl_0_225 br_0_225 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c225
*+ bl_0_225 br_0_225 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c225
*+ bl_0_225 br_0_225 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c225
*+ bl_0_225 br_0_225 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c225
*+ bl_0_225 br_0_225 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c225
*+ bl_0_225 br_0_225 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c225
*+ bl_0_225 br_0_225 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c225
*+ bl_0_225 br_0_225 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c225
*+ bl_0_225 br_0_225 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c225
*+ bl_0_225 br_0_225 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c225
*+ bl_0_225 br_0_225 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c225
*+ bl_0_225 br_0_225 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c225
*+ bl_0_225 br_0_225 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c225
*+ bl_0_225 br_0_225 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c225
*+ bl_0_225 br_0_225 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c225
*+ bl_0_225 br_0_225 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c225
*+ bl_0_225 br_0_225 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c225
*+ bl_0_225 br_0_225 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c225
*+ bl_0_225 br_0_225 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c225
*+ bl_0_225 br_0_225 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c225
*+ bl_0_225 br_0_225 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c225
*+ bl_0_225 br_0_225 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c225
*+ bl_0_225 br_0_225 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c225
*+ bl_0_225 br_0_225 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c225
*+ bl_0_225 br_0_225 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c225
*+ bl_0_225 br_0_225 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c225
*+ bl_0_225 br_0_225 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c225
*+ bl_0_225 br_0_225 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c225
*+ bl_0_225 br_0_225 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c225
*+ bl_0_225 br_0_225 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c225
*+ bl_0_225 br_0_225 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c225
*+ bl_0_225 br_0_225 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c225
*+ bl_0_225 br_0_225 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c225
*+ bl_0_225 br_0_225 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c225
*+ bl_0_225 br_0_225 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c225
*+ bl_0_225 br_0_225 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c225
*+ bl_0_225 br_0_225 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c225
*+ bl_0_225 br_0_225 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c225
*+ bl_0_225 br_0_225 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c225
*+ bl_0_225 br_0_225 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c225
*+ bl_0_225 br_0_225 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c225
*+ bl_0_225 br_0_225 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c225
*+ bl_0_225 br_0_225 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c225
*+ bl_0_225 br_0_225 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c225
*+ bl_0_225 br_0_225 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c225
*+ bl_0_225 br_0_225 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c225
*+ bl_0_225 br_0_225 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c225
*+ bl_0_225 br_0_225 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c225
*+ bl_0_225 br_0_225 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c225
*+ bl_0_225 br_0_225 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c225
*+ bl_0_225 br_0_225 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c225
*+ bl_0_225 br_0_225 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c225
*+ bl_0_225 br_0_225 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c225
*+ bl_0_225 br_0_225 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c225
*+ bl_0_225 br_0_225 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c225
*+ bl_0_225 br_0_225 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c225
*+ bl_0_225 br_0_225 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c225
*+ bl_0_225 br_0_225 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c225
*+ bl_0_225 br_0_225 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c225
*+ bl_0_225 br_0_225 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c225
*+ bl_0_225 br_0_225 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c225
*+ bl_0_225 br_0_225 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c225
*+ bl_0_225 br_0_225 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c225
*+ bl_0_225 br_0_225 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c225
*+ bl_0_225 br_0_225 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c225
*+ bl_0_225 br_0_225 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c225
*+ bl_0_225 br_0_225 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c225
*+ bl_0_225 br_0_225 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c225
*+ bl_0_225 br_0_225 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c225
*+ bl_0_225 br_0_225 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c225
*+ bl_0_225 br_0_225 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c225
*+ bl_0_225 br_0_225 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c225
*+ bl_0_225 br_0_225 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c225
*+ bl_0_225 br_0_225 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c225
*+ bl_0_225 br_0_225 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c225
*+ bl_0_225 br_0_225 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c225
*+ bl_0_225 br_0_225 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c225
*+ bl_0_225 br_0_225 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c225
+ bl_0_225 br_0_225 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c226
+ bl_0_226 br_0_226 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c226
*+ bl_0_226 br_0_226 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c226
*+ bl_0_226 br_0_226 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c226
*+ bl_0_226 br_0_226 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c226
*+ bl_0_226 br_0_226 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c226
*+ bl_0_226 br_0_226 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c226
*+ bl_0_226 br_0_226 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c226
*+ bl_0_226 br_0_226 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c226
*+ bl_0_226 br_0_226 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c226
*+ bl_0_226 br_0_226 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c226
*+ bl_0_226 br_0_226 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c226
*+ bl_0_226 br_0_226 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c226
*+ bl_0_226 br_0_226 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c226
*+ bl_0_226 br_0_226 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c226
*+ bl_0_226 br_0_226 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c226
*+ bl_0_226 br_0_226 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c226
*+ bl_0_226 br_0_226 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c226
*+ bl_0_226 br_0_226 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c226
*+ bl_0_226 br_0_226 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c226
*+ bl_0_226 br_0_226 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c226
*+ bl_0_226 br_0_226 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c226
*+ bl_0_226 br_0_226 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c226
*+ bl_0_226 br_0_226 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c226
*+ bl_0_226 br_0_226 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c226
*+ bl_0_226 br_0_226 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c226
*+ bl_0_226 br_0_226 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c226
*+ bl_0_226 br_0_226 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c226
*+ bl_0_226 br_0_226 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c226
*+ bl_0_226 br_0_226 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c226
*+ bl_0_226 br_0_226 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c226
*+ bl_0_226 br_0_226 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c226
*+ bl_0_226 br_0_226 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c226
*+ bl_0_226 br_0_226 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c226
*+ bl_0_226 br_0_226 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c226
*+ bl_0_226 br_0_226 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c226
*+ bl_0_226 br_0_226 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c226
*+ bl_0_226 br_0_226 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c226
*+ bl_0_226 br_0_226 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c226
*+ bl_0_226 br_0_226 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c226
*+ bl_0_226 br_0_226 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c226
*+ bl_0_226 br_0_226 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c226
*+ bl_0_226 br_0_226 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c226
*+ bl_0_226 br_0_226 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c226
*+ bl_0_226 br_0_226 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c226
*+ bl_0_226 br_0_226 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c226
*+ bl_0_226 br_0_226 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c226
*+ bl_0_226 br_0_226 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c226
*+ bl_0_226 br_0_226 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c226
*+ bl_0_226 br_0_226 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c226
*+ bl_0_226 br_0_226 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c226
*+ bl_0_226 br_0_226 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c226
*+ bl_0_226 br_0_226 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c226
*+ bl_0_226 br_0_226 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c226
*+ bl_0_226 br_0_226 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c226
*+ bl_0_226 br_0_226 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c226
*+ bl_0_226 br_0_226 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c226
*+ bl_0_226 br_0_226 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c226
*+ bl_0_226 br_0_226 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c226
*+ bl_0_226 br_0_226 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c226
*+ bl_0_226 br_0_226 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c226
*+ bl_0_226 br_0_226 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c226
*+ bl_0_226 br_0_226 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c226
*+ bl_0_226 br_0_226 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c226
*+ bl_0_226 br_0_226 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c226
*+ bl_0_226 br_0_226 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c226
*+ bl_0_226 br_0_226 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c226
*+ bl_0_226 br_0_226 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c226
*+ bl_0_226 br_0_226 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c226
*+ bl_0_226 br_0_226 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c226
*+ bl_0_226 br_0_226 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c226
*+ bl_0_226 br_0_226 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c226
*+ bl_0_226 br_0_226 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c226
*+ bl_0_226 br_0_226 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c226
*+ bl_0_226 br_0_226 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c226
*+ bl_0_226 br_0_226 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c226
*+ bl_0_226 br_0_226 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c226
*+ bl_0_226 br_0_226 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c226
*+ bl_0_226 br_0_226 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c226
*+ bl_0_226 br_0_226 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c226
*+ bl_0_226 br_0_226 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c226
*+ bl_0_226 br_0_226 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c226
*+ bl_0_226 br_0_226 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c226
*+ bl_0_226 br_0_226 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c226
*+ bl_0_226 br_0_226 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c226
*+ bl_0_226 br_0_226 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c226
*+ bl_0_226 br_0_226 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c226
*+ bl_0_226 br_0_226 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c226
*+ bl_0_226 br_0_226 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c226
*+ bl_0_226 br_0_226 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c226
*+ bl_0_226 br_0_226 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c226
*+ bl_0_226 br_0_226 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c226
*+ bl_0_226 br_0_226 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c226
*+ bl_0_226 br_0_226 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c226
*+ bl_0_226 br_0_226 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c226
*+ bl_0_226 br_0_226 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c226
*+ bl_0_226 br_0_226 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c226
*+ bl_0_226 br_0_226 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c226
*+ bl_0_226 br_0_226 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c226
*+ bl_0_226 br_0_226 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c226
*+ bl_0_226 br_0_226 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c226
*+ bl_0_226 br_0_226 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c226
*+ bl_0_226 br_0_226 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c226
*+ bl_0_226 br_0_226 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c226
*+ bl_0_226 br_0_226 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c226
*+ bl_0_226 br_0_226 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c226
*+ bl_0_226 br_0_226 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c226
*+ bl_0_226 br_0_226 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c226
*+ bl_0_226 br_0_226 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c226
*+ bl_0_226 br_0_226 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c226
*+ bl_0_226 br_0_226 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c226
*+ bl_0_226 br_0_226 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c226
*+ bl_0_226 br_0_226 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c226
*+ bl_0_226 br_0_226 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c226
*+ bl_0_226 br_0_226 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c226
*+ bl_0_226 br_0_226 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c226
*+ bl_0_226 br_0_226 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c226
*+ bl_0_226 br_0_226 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c226
*+ bl_0_226 br_0_226 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c226
*+ bl_0_226 br_0_226 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c226
*+ bl_0_226 br_0_226 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c226
*+ bl_0_226 br_0_226 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c226
*+ bl_0_226 br_0_226 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c226
*+ bl_0_226 br_0_226 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c226
*+ bl_0_226 br_0_226 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c226
*+ bl_0_226 br_0_226 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c226
*+ bl_0_226 br_0_226 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c226
*+ bl_0_226 br_0_226 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c226
+ bl_0_226 br_0_226 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c227
+ bl_0_227 br_0_227 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c227
*+ bl_0_227 br_0_227 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c227
*+ bl_0_227 br_0_227 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c227
*+ bl_0_227 br_0_227 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c227
*+ bl_0_227 br_0_227 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c227
*+ bl_0_227 br_0_227 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c227
*+ bl_0_227 br_0_227 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c227
*+ bl_0_227 br_0_227 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c227
*+ bl_0_227 br_0_227 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c227
*+ bl_0_227 br_0_227 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c227
*+ bl_0_227 br_0_227 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c227
*+ bl_0_227 br_0_227 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c227
*+ bl_0_227 br_0_227 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c227
*+ bl_0_227 br_0_227 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c227
*+ bl_0_227 br_0_227 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c227
*+ bl_0_227 br_0_227 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c227
*+ bl_0_227 br_0_227 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c227
*+ bl_0_227 br_0_227 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c227
*+ bl_0_227 br_0_227 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c227
*+ bl_0_227 br_0_227 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c227
*+ bl_0_227 br_0_227 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c227
*+ bl_0_227 br_0_227 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c227
*+ bl_0_227 br_0_227 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c227
*+ bl_0_227 br_0_227 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c227
*+ bl_0_227 br_0_227 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c227
*+ bl_0_227 br_0_227 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c227
*+ bl_0_227 br_0_227 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c227
*+ bl_0_227 br_0_227 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c227
*+ bl_0_227 br_0_227 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c227
*+ bl_0_227 br_0_227 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c227
*+ bl_0_227 br_0_227 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c227
*+ bl_0_227 br_0_227 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c227
*+ bl_0_227 br_0_227 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c227
*+ bl_0_227 br_0_227 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c227
*+ bl_0_227 br_0_227 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c227
*+ bl_0_227 br_0_227 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c227
*+ bl_0_227 br_0_227 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c227
*+ bl_0_227 br_0_227 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c227
*+ bl_0_227 br_0_227 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c227
*+ bl_0_227 br_0_227 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c227
*+ bl_0_227 br_0_227 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c227
*+ bl_0_227 br_0_227 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c227
*+ bl_0_227 br_0_227 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c227
*+ bl_0_227 br_0_227 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c227
*+ bl_0_227 br_0_227 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c227
*+ bl_0_227 br_0_227 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c227
*+ bl_0_227 br_0_227 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c227
*+ bl_0_227 br_0_227 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c227
*+ bl_0_227 br_0_227 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c227
*+ bl_0_227 br_0_227 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c227
*+ bl_0_227 br_0_227 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c227
*+ bl_0_227 br_0_227 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c227
*+ bl_0_227 br_0_227 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c227
*+ bl_0_227 br_0_227 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c227
*+ bl_0_227 br_0_227 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c227
*+ bl_0_227 br_0_227 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c227
*+ bl_0_227 br_0_227 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c227
*+ bl_0_227 br_0_227 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c227
*+ bl_0_227 br_0_227 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c227
*+ bl_0_227 br_0_227 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c227
*+ bl_0_227 br_0_227 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c227
*+ bl_0_227 br_0_227 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c227
*+ bl_0_227 br_0_227 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c227
*+ bl_0_227 br_0_227 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c227
*+ bl_0_227 br_0_227 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c227
*+ bl_0_227 br_0_227 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c227
*+ bl_0_227 br_0_227 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c227
*+ bl_0_227 br_0_227 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c227
*+ bl_0_227 br_0_227 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c227
*+ bl_0_227 br_0_227 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c227
*+ bl_0_227 br_0_227 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c227
*+ bl_0_227 br_0_227 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c227
*+ bl_0_227 br_0_227 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c227
*+ bl_0_227 br_0_227 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c227
*+ bl_0_227 br_0_227 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c227
*+ bl_0_227 br_0_227 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c227
*+ bl_0_227 br_0_227 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c227
*+ bl_0_227 br_0_227 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c227
*+ bl_0_227 br_0_227 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c227
*+ bl_0_227 br_0_227 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c227
*+ bl_0_227 br_0_227 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c227
*+ bl_0_227 br_0_227 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c227
*+ bl_0_227 br_0_227 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c227
*+ bl_0_227 br_0_227 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c227
*+ bl_0_227 br_0_227 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c227
*+ bl_0_227 br_0_227 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c227
*+ bl_0_227 br_0_227 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c227
*+ bl_0_227 br_0_227 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c227
*+ bl_0_227 br_0_227 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c227
*+ bl_0_227 br_0_227 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c227
*+ bl_0_227 br_0_227 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c227
*+ bl_0_227 br_0_227 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c227
*+ bl_0_227 br_0_227 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c227
*+ bl_0_227 br_0_227 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c227
*+ bl_0_227 br_0_227 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c227
*+ bl_0_227 br_0_227 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c227
*+ bl_0_227 br_0_227 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c227
*+ bl_0_227 br_0_227 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c227
*+ bl_0_227 br_0_227 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c227
*+ bl_0_227 br_0_227 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c227
*+ bl_0_227 br_0_227 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c227
*+ bl_0_227 br_0_227 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c227
*+ bl_0_227 br_0_227 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c227
*+ bl_0_227 br_0_227 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c227
*+ bl_0_227 br_0_227 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c227
*+ bl_0_227 br_0_227 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c227
*+ bl_0_227 br_0_227 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c227
*+ bl_0_227 br_0_227 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c227
*+ bl_0_227 br_0_227 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c227
*+ bl_0_227 br_0_227 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c227
*+ bl_0_227 br_0_227 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c227
*+ bl_0_227 br_0_227 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c227
*+ bl_0_227 br_0_227 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c227
*+ bl_0_227 br_0_227 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c227
*+ bl_0_227 br_0_227 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c227
*+ bl_0_227 br_0_227 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c227
*+ bl_0_227 br_0_227 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c227
*+ bl_0_227 br_0_227 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c227
*+ bl_0_227 br_0_227 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c227
*+ bl_0_227 br_0_227 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c227
*+ bl_0_227 br_0_227 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c227
*+ bl_0_227 br_0_227 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c227
*+ bl_0_227 br_0_227 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c227
*+ bl_0_227 br_0_227 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c227
*+ bl_0_227 br_0_227 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c227
*+ bl_0_227 br_0_227 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c227
*+ bl_0_227 br_0_227 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c227
+ bl_0_227 br_0_227 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c228
+ bl_0_228 br_0_228 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c228
*+ bl_0_228 br_0_228 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c228
*+ bl_0_228 br_0_228 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c228
*+ bl_0_228 br_0_228 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c228
*+ bl_0_228 br_0_228 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c228
*+ bl_0_228 br_0_228 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c228
*+ bl_0_228 br_0_228 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c228
*+ bl_0_228 br_0_228 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c228
*+ bl_0_228 br_0_228 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c228
*+ bl_0_228 br_0_228 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c228
*+ bl_0_228 br_0_228 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c228
*+ bl_0_228 br_0_228 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c228
*+ bl_0_228 br_0_228 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c228
*+ bl_0_228 br_0_228 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c228
*+ bl_0_228 br_0_228 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c228
*+ bl_0_228 br_0_228 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c228
*+ bl_0_228 br_0_228 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c228
*+ bl_0_228 br_0_228 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c228
*+ bl_0_228 br_0_228 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c228
*+ bl_0_228 br_0_228 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c228
*+ bl_0_228 br_0_228 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c228
*+ bl_0_228 br_0_228 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c228
*+ bl_0_228 br_0_228 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c228
*+ bl_0_228 br_0_228 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c228
*+ bl_0_228 br_0_228 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c228
*+ bl_0_228 br_0_228 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c228
*+ bl_0_228 br_0_228 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c228
*+ bl_0_228 br_0_228 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c228
*+ bl_0_228 br_0_228 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c228
*+ bl_0_228 br_0_228 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c228
*+ bl_0_228 br_0_228 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c228
*+ bl_0_228 br_0_228 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c228
*+ bl_0_228 br_0_228 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c228
*+ bl_0_228 br_0_228 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c228
*+ bl_0_228 br_0_228 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c228
*+ bl_0_228 br_0_228 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c228
*+ bl_0_228 br_0_228 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c228
*+ bl_0_228 br_0_228 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c228
*+ bl_0_228 br_0_228 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c228
*+ bl_0_228 br_0_228 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c228
*+ bl_0_228 br_0_228 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c228
*+ bl_0_228 br_0_228 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c228
*+ bl_0_228 br_0_228 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c228
*+ bl_0_228 br_0_228 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c228
*+ bl_0_228 br_0_228 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c228
*+ bl_0_228 br_0_228 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c228
*+ bl_0_228 br_0_228 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c228
*+ bl_0_228 br_0_228 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c228
*+ bl_0_228 br_0_228 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c228
*+ bl_0_228 br_0_228 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c228
*+ bl_0_228 br_0_228 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c228
*+ bl_0_228 br_0_228 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c228
*+ bl_0_228 br_0_228 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c228
*+ bl_0_228 br_0_228 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c228
*+ bl_0_228 br_0_228 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c228
*+ bl_0_228 br_0_228 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c228
*+ bl_0_228 br_0_228 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c228
*+ bl_0_228 br_0_228 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c228
*+ bl_0_228 br_0_228 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c228
*+ bl_0_228 br_0_228 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c228
*+ bl_0_228 br_0_228 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c228
*+ bl_0_228 br_0_228 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c228
*+ bl_0_228 br_0_228 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c228
*+ bl_0_228 br_0_228 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c228
*+ bl_0_228 br_0_228 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c228
*+ bl_0_228 br_0_228 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c228
*+ bl_0_228 br_0_228 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c228
*+ bl_0_228 br_0_228 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c228
*+ bl_0_228 br_0_228 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c228
*+ bl_0_228 br_0_228 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c228
*+ bl_0_228 br_0_228 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c228
*+ bl_0_228 br_0_228 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c228
*+ bl_0_228 br_0_228 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c228
*+ bl_0_228 br_0_228 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c228
*+ bl_0_228 br_0_228 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c228
*+ bl_0_228 br_0_228 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c228
*+ bl_0_228 br_0_228 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c228
*+ bl_0_228 br_0_228 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c228
*+ bl_0_228 br_0_228 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c228
*+ bl_0_228 br_0_228 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c228
*+ bl_0_228 br_0_228 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c228
*+ bl_0_228 br_0_228 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c228
*+ bl_0_228 br_0_228 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c228
*+ bl_0_228 br_0_228 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c228
*+ bl_0_228 br_0_228 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c228
*+ bl_0_228 br_0_228 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c228
*+ bl_0_228 br_0_228 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c228
*+ bl_0_228 br_0_228 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c228
*+ bl_0_228 br_0_228 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c228
*+ bl_0_228 br_0_228 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c228
*+ bl_0_228 br_0_228 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c228
*+ bl_0_228 br_0_228 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c228
*+ bl_0_228 br_0_228 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c228
*+ bl_0_228 br_0_228 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c228
*+ bl_0_228 br_0_228 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c228
*+ bl_0_228 br_0_228 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c228
*+ bl_0_228 br_0_228 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c228
*+ bl_0_228 br_0_228 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c228
*+ bl_0_228 br_0_228 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c228
*+ bl_0_228 br_0_228 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c228
*+ bl_0_228 br_0_228 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c228
*+ bl_0_228 br_0_228 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c228
*+ bl_0_228 br_0_228 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c228
*+ bl_0_228 br_0_228 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c228
*+ bl_0_228 br_0_228 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c228
*+ bl_0_228 br_0_228 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c228
*+ bl_0_228 br_0_228 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c228
*+ bl_0_228 br_0_228 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c228
*+ bl_0_228 br_0_228 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c228
*+ bl_0_228 br_0_228 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c228
*+ bl_0_228 br_0_228 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c228
*+ bl_0_228 br_0_228 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c228
*+ bl_0_228 br_0_228 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c228
*+ bl_0_228 br_0_228 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c228
*+ bl_0_228 br_0_228 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c228
*+ bl_0_228 br_0_228 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c228
*+ bl_0_228 br_0_228 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c228
*+ bl_0_228 br_0_228 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c228
*+ bl_0_228 br_0_228 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c228
*+ bl_0_228 br_0_228 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c228
*+ bl_0_228 br_0_228 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c228
*+ bl_0_228 br_0_228 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c228
*+ bl_0_228 br_0_228 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c228
*+ bl_0_228 br_0_228 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c228
*+ bl_0_228 br_0_228 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c228
*+ bl_0_228 br_0_228 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c228
*+ bl_0_228 br_0_228 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c228
+ bl_0_228 br_0_228 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c229
+ bl_0_229 br_0_229 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c229
*+ bl_0_229 br_0_229 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c229
*+ bl_0_229 br_0_229 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c229
*+ bl_0_229 br_0_229 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c229
*+ bl_0_229 br_0_229 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c229
*+ bl_0_229 br_0_229 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c229
*+ bl_0_229 br_0_229 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c229
*+ bl_0_229 br_0_229 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c229
*+ bl_0_229 br_0_229 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c229
*+ bl_0_229 br_0_229 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c229
*+ bl_0_229 br_0_229 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c229
*+ bl_0_229 br_0_229 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c229
*+ bl_0_229 br_0_229 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c229
*+ bl_0_229 br_0_229 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c229
*+ bl_0_229 br_0_229 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c229
*+ bl_0_229 br_0_229 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c229
*+ bl_0_229 br_0_229 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c229
*+ bl_0_229 br_0_229 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c229
*+ bl_0_229 br_0_229 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c229
*+ bl_0_229 br_0_229 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c229
*+ bl_0_229 br_0_229 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c229
*+ bl_0_229 br_0_229 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c229
*+ bl_0_229 br_0_229 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c229
*+ bl_0_229 br_0_229 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c229
*+ bl_0_229 br_0_229 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c229
*+ bl_0_229 br_0_229 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c229
*+ bl_0_229 br_0_229 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c229
*+ bl_0_229 br_0_229 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c229
*+ bl_0_229 br_0_229 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c229
*+ bl_0_229 br_0_229 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c229
*+ bl_0_229 br_0_229 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c229
*+ bl_0_229 br_0_229 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c229
*+ bl_0_229 br_0_229 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c229
*+ bl_0_229 br_0_229 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c229
*+ bl_0_229 br_0_229 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c229
*+ bl_0_229 br_0_229 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c229
*+ bl_0_229 br_0_229 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c229
*+ bl_0_229 br_0_229 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c229
*+ bl_0_229 br_0_229 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c229
*+ bl_0_229 br_0_229 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c229
*+ bl_0_229 br_0_229 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c229
*+ bl_0_229 br_0_229 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c229
*+ bl_0_229 br_0_229 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c229
*+ bl_0_229 br_0_229 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c229
*+ bl_0_229 br_0_229 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c229
*+ bl_0_229 br_0_229 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c229
*+ bl_0_229 br_0_229 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c229
*+ bl_0_229 br_0_229 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c229
*+ bl_0_229 br_0_229 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c229
*+ bl_0_229 br_0_229 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c229
*+ bl_0_229 br_0_229 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c229
*+ bl_0_229 br_0_229 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c229
*+ bl_0_229 br_0_229 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c229
*+ bl_0_229 br_0_229 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c229
*+ bl_0_229 br_0_229 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c229
*+ bl_0_229 br_0_229 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c229
*+ bl_0_229 br_0_229 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c229
*+ bl_0_229 br_0_229 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c229
*+ bl_0_229 br_0_229 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c229
*+ bl_0_229 br_0_229 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c229
*+ bl_0_229 br_0_229 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c229
*+ bl_0_229 br_0_229 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c229
*+ bl_0_229 br_0_229 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c229
*+ bl_0_229 br_0_229 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c229
*+ bl_0_229 br_0_229 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c229
*+ bl_0_229 br_0_229 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c229
*+ bl_0_229 br_0_229 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c229
*+ bl_0_229 br_0_229 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c229
*+ bl_0_229 br_0_229 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c229
*+ bl_0_229 br_0_229 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c229
*+ bl_0_229 br_0_229 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c229
*+ bl_0_229 br_0_229 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c229
*+ bl_0_229 br_0_229 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c229
*+ bl_0_229 br_0_229 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c229
*+ bl_0_229 br_0_229 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c229
*+ bl_0_229 br_0_229 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c229
*+ bl_0_229 br_0_229 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c229
*+ bl_0_229 br_0_229 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c229
*+ bl_0_229 br_0_229 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c229
*+ bl_0_229 br_0_229 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c229
*+ bl_0_229 br_0_229 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c229
*+ bl_0_229 br_0_229 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c229
*+ bl_0_229 br_0_229 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c229
*+ bl_0_229 br_0_229 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c229
*+ bl_0_229 br_0_229 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c229
*+ bl_0_229 br_0_229 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c229
*+ bl_0_229 br_0_229 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c229
*+ bl_0_229 br_0_229 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c229
*+ bl_0_229 br_0_229 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c229
*+ bl_0_229 br_0_229 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c229
*+ bl_0_229 br_0_229 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c229
*+ bl_0_229 br_0_229 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c229
*+ bl_0_229 br_0_229 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c229
*+ bl_0_229 br_0_229 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c229
*+ bl_0_229 br_0_229 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c229
*+ bl_0_229 br_0_229 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c229
*+ bl_0_229 br_0_229 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c229
*+ bl_0_229 br_0_229 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c229
*+ bl_0_229 br_0_229 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c229
*+ bl_0_229 br_0_229 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c229
*+ bl_0_229 br_0_229 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c229
*+ bl_0_229 br_0_229 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c229
*+ bl_0_229 br_0_229 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c229
*+ bl_0_229 br_0_229 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c229
*+ bl_0_229 br_0_229 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c229
*+ bl_0_229 br_0_229 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c229
*+ bl_0_229 br_0_229 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c229
*+ bl_0_229 br_0_229 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c229
*+ bl_0_229 br_0_229 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c229
*+ bl_0_229 br_0_229 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c229
*+ bl_0_229 br_0_229 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c229
*+ bl_0_229 br_0_229 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c229
*+ bl_0_229 br_0_229 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c229
*+ bl_0_229 br_0_229 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c229
*+ bl_0_229 br_0_229 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c229
*+ bl_0_229 br_0_229 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c229
*+ bl_0_229 br_0_229 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c229
*+ bl_0_229 br_0_229 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c229
*+ bl_0_229 br_0_229 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c229
*+ bl_0_229 br_0_229 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c229
*+ bl_0_229 br_0_229 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c229
*+ bl_0_229 br_0_229 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c229
*+ bl_0_229 br_0_229 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c229
*+ bl_0_229 br_0_229 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c229
*+ bl_0_229 br_0_229 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c229
*+ bl_0_229 br_0_229 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c229
*+ bl_0_229 br_0_229 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c229
+ bl_0_229 br_0_229 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c230
+ bl_0_230 br_0_230 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c230
*+ bl_0_230 br_0_230 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c230
*+ bl_0_230 br_0_230 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c230
*+ bl_0_230 br_0_230 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c230
*+ bl_0_230 br_0_230 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c230
*+ bl_0_230 br_0_230 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c230
*+ bl_0_230 br_0_230 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c230
*+ bl_0_230 br_0_230 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c230
*+ bl_0_230 br_0_230 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c230
*+ bl_0_230 br_0_230 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c230
*+ bl_0_230 br_0_230 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c230
*+ bl_0_230 br_0_230 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c230
*+ bl_0_230 br_0_230 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c230
*+ bl_0_230 br_0_230 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c230
*+ bl_0_230 br_0_230 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c230
*+ bl_0_230 br_0_230 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c230
*+ bl_0_230 br_0_230 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c230
*+ bl_0_230 br_0_230 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c230
*+ bl_0_230 br_0_230 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c230
*+ bl_0_230 br_0_230 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c230
*+ bl_0_230 br_0_230 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c230
*+ bl_0_230 br_0_230 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c230
*+ bl_0_230 br_0_230 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c230
*+ bl_0_230 br_0_230 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c230
*+ bl_0_230 br_0_230 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c230
*+ bl_0_230 br_0_230 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c230
*+ bl_0_230 br_0_230 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c230
*+ bl_0_230 br_0_230 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c230
*+ bl_0_230 br_0_230 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c230
*+ bl_0_230 br_0_230 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c230
*+ bl_0_230 br_0_230 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c230
*+ bl_0_230 br_0_230 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c230
*+ bl_0_230 br_0_230 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c230
*+ bl_0_230 br_0_230 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c230
*+ bl_0_230 br_0_230 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c230
*+ bl_0_230 br_0_230 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c230
*+ bl_0_230 br_0_230 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c230
*+ bl_0_230 br_0_230 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c230
*+ bl_0_230 br_0_230 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c230
*+ bl_0_230 br_0_230 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c230
*+ bl_0_230 br_0_230 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c230
*+ bl_0_230 br_0_230 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c230
*+ bl_0_230 br_0_230 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c230
*+ bl_0_230 br_0_230 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c230
*+ bl_0_230 br_0_230 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c230
*+ bl_0_230 br_0_230 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c230
*+ bl_0_230 br_0_230 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c230
*+ bl_0_230 br_0_230 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c230
*+ bl_0_230 br_0_230 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c230
*+ bl_0_230 br_0_230 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c230
*+ bl_0_230 br_0_230 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c230
*+ bl_0_230 br_0_230 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c230
*+ bl_0_230 br_0_230 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c230
*+ bl_0_230 br_0_230 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c230
*+ bl_0_230 br_0_230 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c230
*+ bl_0_230 br_0_230 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c230
*+ bl_0_230 br_0_230 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c230
*+ bl_0_230 br_0_230 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c230
*+ bl_0_230 br_0_230 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c230
*+ bl_0_230 br_0_230 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c230
*+ bl_0_230 br_0_230 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c230
*+ bl_0_230 br_0_230 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c230
*+ bl_0_230 br_0_230 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c230
*+ bl_0_230 br_0_230 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c230
*+ bl_0_230 br_0_230 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c230
*+ bl_0_230 br_0_230 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c230
*+ bl_0_230 br_0_230 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c230
*+ bl_0_230 br_0_230 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c230
*+ bl_0_230 br_0_230 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c230
*+ bl_0_230 br_0_230 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c230
*+ bl_0_230 br_0_230 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c230
*+ bl_0_230 br_0_230 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c230
*+ bl_0_230 br_0_230 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c230
*+ bl_0_230 br_0_230 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c230
*+ bl_0_230 br_0_230 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c230
*+ bl_0_230 br_0_230 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c230
*+ bl_0_230 br_0_230 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c230
*+ bl_0_230 br_0_230 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c230
*+ bl_0_230 br_0_230 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c230
*+ bl_0_230 br_0_230 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c230
*+ bl_0_230 br_0_230 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c230
*+ bl_0_230 br_0_230 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c230
*+ bl_0_230 br_0_230 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c230
*+ bl_0_230 br_0_230 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c230
*+ bl_0_230 br_0_230 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c230
*+ bl_0_230 br_0_230 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c230
*+ bl_0_230 br_0_230 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c230
*+ bl_0_230 br_0_230 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c230
*+ bl_0_230 br_0_230 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c230
*+ bl_0_230 br_0_230 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c230
*+ bl_0_230 br_0_230 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c230
*+ bl_0_230 br_0_230 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c230
*+ bl_0_230 br_0_230 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c230
*+ bl_0_230 br_0_230 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c230
*+ bl_0_230 br_0_230 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c230
*+ bl_0_230 br_0_230 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c230
*+ bl_0_230 br_0_230 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c230
*+ bl_0_230 br_0_230 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c230
*+ bl_0_230 br_0_230 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c230
*+ bl_0_230 br_0_230 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c230
*+ bl_0_230 br_0_230 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c230
*+ bl_0_230 br_0_230 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c230
*+ bl_0_230 br_0_230 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c230
*+ bl_0_230 br_0_230 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c230
*+ bl_0_230 br_0_230 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c230
*+ bl_0_230 br_0_230 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c230
*+ bl_0_230 br_0_230 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c230
*+ bl_0_230 br_0_230 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c230
*+ bl_0_230 br_0_230 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c230
*+ bl_0_230 br_0_230 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c230
*+ bl_0_230 br_0_230 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c230
*+ bl_0_230 br_0_230 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c230
*+ bl_0_230 br_0_230 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c230
*+ bl_0_230 br_0_230 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c230
*+ bl_0_230 br_0_230 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c230
*+ bl_0_230 br_0_230 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c230
*+ bl_0_230 br_0_230 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c230
*+ bl_0_230 br_0_230 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c230
*+ bl_0_230 br_0_230 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c230
*+ bl_0_230 br_0_230 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c230
*+ bl_0_230 br_0_230 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c230
*+ bl_0_230 br_0_230 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c230
*+ bl_0_230 br_0_230 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c230
*+ bl_0_230 br_0_230 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c230
*+ bl_0_230 br_0_230 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c230
*+ bl_0_230 br_0_230 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c230
*+ bl_0_230 br_0_230 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c230
+ bl_0_230 br_0_230 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c231
+ bl_0_231 br_0_231 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c231
*+ bl_0_231 br_0_231 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c231
*+ bl_0_231 br_0_231 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c231
*+ bl_0_231 br_0_231 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c231
*+ bl_0_231 br_0_231 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c231
*+ bl_0_231 br_0_231 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c231
*+ bl_0_231 br_0_231 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c231
*+ bl_0_231 br_0_231 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c231
*+ bl_0_231 br_0_231 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c231
*+ bl_0_231 br_0_231 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c231
*+ bl_0_231 br_0_231 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c231
*+ bl_0_231 br_0_231 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c231
*+ bl_0_231 br_0_231 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c231
*+ bl_0_231 br_0_231 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c231
*+ bl_0_231 br_0_231 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c231
*+ bl_0_231 br_0_231 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c231
*+ bl_0_231 br_0_231 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c231
*+ bl_0_231 br_0_231 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c231
*+ bl_0_231 br_0_231 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c231
*+ bl_0_231 br_0_231 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c231
*+ bl_0_231 br_0_231 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c231
*+ bl_0_231 br_0_231 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c231
*+ bl_0_231 br_0_231 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c231
*+ bl_0_231 br_0_231 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c231
*+ bl_0_231 br_0_231 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c231
*+ bl_0_231 br_0_231 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c231
*+ bl_0_231 br_0_231 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c231
*+ bl_0_231 br_0_231 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c231
*+ bl_0_231 br_0_231 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c231
*+ bl_0_231 br_0_231 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c231
*+ bl_0_231 br_0_231 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c231
*+ bl_0_231 br_0_231 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c231
*+ bl_0_231 br_0_231 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c231
*+ bl_0_231 br_0_231 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c231
*+ bl_0_231 br_0_231 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c231
*+ bl_0_231 br_0_231 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c231
*+ bl_0_231 br_0_231 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c231
*+ bl_0_231 br_0_231 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c231
*+ bl_0_231 br_0_231 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c231
*+ bl_0_231 br_0_231 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c231
*+ bl_0_231 br_0_231 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c231
*+ bl_0_231 br_0_231 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c231
*+ bl_0_231 br_0_231 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c231
*+ bl_0_231 br_0_231 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c231
*+ bl_0_231 br_0_231 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c231
*+ bl_0_231 br_0_231 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c231
*+ bl_0_231 br_0_231 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c231
*+ bl_0_231 br_0_231 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c231
*+ bl_0_231 br_0_231 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c231
*+ bl_0_231 br_0_231 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c231
*+ bl_0_231 br_0_231 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c231
*+ bl_0_231 br_0_231 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c231
*+ bl_0_231 br_0_231 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c231
*+ bl_0_231 br_0_231 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c231
*+ bl_0_231 br_0_231 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c231
*+ bl_0_231 br_0_231 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c231
*+ bl_0_231 br_0_231 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c231
*+ bl_0_231 br_0_231 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c231
*+ bl_0_231 br_0_231 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c231
*+ bl_0_231 br_0_231 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c231
*+ bl_0_231 br_0_231 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c231
*+ bl_0_231 br_0_231 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c231
*+ bl_0_231 br_0_231 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c231
*+ bl_0_231 br_0_231 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c231
*+ bl_0_231 br_0_231 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c231
*+ bl_0_231 br_0_231 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c231
*+ bl_0_231 br_0_231 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c231
*+ bl_0_231 br_0_231 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c231
*+ bl_0_231 br_0_231 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c231
*+ bl_0_231 br_0_231 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c231
*+ bl_0_231 br_0_231 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c231
*+ bl_0_231 br_0_231 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c231
*+ bl_0_231 br_0_231 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c231
*+ bl_0_231 br_0_231 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c231
*+ bl_0_231 br_0_231 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c231
*+ bl_0_231 br_0_231 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c231
*+ bl_0_231 br_0_231 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c231
*+ bl_0_231 br_0_231 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c231
*+ bl_0_231 br_0_231 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c231
*+ bl_0_231 br_0_231 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c231
*+ bl_0_231 br_0_231 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c231
*+ bl_0_231 br_0_231 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c231
*+ bl_0_231 br_0_231 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c231
*+ bl_0_231 br_0_231 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c231
*+ bl_0_231 br_0_231 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c231
*+ bl_0_231 br_0_231 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c231
*+ bl_0_231 br_0_231 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c231
*+ bl_0_231 br_0_231 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c231
*+ bl_0_231 br_0_231 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c231
*+ bl_0_231 br_0_231 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c231
*+ bl_0_231 br_0_231 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c231
*+ bl_0_231 br_0_231 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c231
*+ bl_0_231 br_0_231 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c231
*+ bl_0_231 br_0_231 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c231
*+ bl_0_231 br_0_231 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c231
*+ bl_0_231 br_0_231 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c231
*+ bl_0_231 br_0_231 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c231
*+ bl_0_231 br_0_231 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c231
*+ bl_0_231 br_0_231 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c231
*+ bl_0_231 br_0_231 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c231
*+ bl_0_231 br_0_231 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c231
*+ bl_0_231 br_0_231 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c231
*+ bl_0_231 br_0_231 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c231
*+ bl_0_231 br_0_231 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c231
*+ bl_0_231 br_0_231 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c231
*+ bl_0_231 br_0_231 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c231
*+ bl_0_231 br_0_231 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c231
*+ bl_0_231 br_0_231 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c231
*+ bl_0_231 br_0_231 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c231
*+ bl_0_231 br_0_231 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c231
*+ bl_0_231 br_0_231 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c231
*+ bl_0_231 br_0_231 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c231
*+ bl_0_231 br_0_231 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c231
*+ bl_0_231 br_0_231 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c231
*+ bl_0_231 br_0_231 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c231
*+ bl_0_231 br_0_231 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c231
*+ bl_0_231 br_0_231 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c231
*+ bl_0_231 br_0_231 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c231
*+ bl_0_231 br_0_231 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c231
*+ bl_0_231 br_0_231 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c231
*+ bl_0_231 br_0_231 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c231
*+ bl_0_231 br_0_231 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c231
*+ bl_0_231 br_0_231 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c231
*+ bl_0_231 br_0_231 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c231
*+ bl_0_231 br_0_231 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c231
*+ bl_0_231 br_0_231 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c231
*+ bl_0_231 br_0_231 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c231
+ bl_0_231 br_0_231 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c232
+ bl_0_232 br_0_232 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c232
*+ bl_0_232 br_0_232 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c232
*+ bl_0_232 br_0_232 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c232
*+ bl_0_232 br_0_232 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c232
*+ bl_0_232 br_0_232 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c232
*+ bl_0_232 br_0_232 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c232
*+ bl_0_232 br_0_232 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c232
*+ bl_0_232 br_0_232 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c232
*+ bl_0_232 br_0_232 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c232
*+ bl_0_232 br_0_232 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c232
*+ bl_0_232 br_0_232 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c232
*+ bl_0_232 br_0_232 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c232
*+ bl_0_232 br_0_232 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c232
*+ bl_0_232 br_0_232 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c232
*+ bl_0_232 br_0_232 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c232
*+ bl_0_232 br_0_232 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c232
*+ bl_0_232 br_0_232 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c232
*+ bl_0_232 br_0_232 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c232
*+ bl_0_232 br_0_232 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c232
*+ bl_0_232 br_0_232 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c232
*+ bl_0_232 br_0_232 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c232
*+ bl_0_232 br_0_232 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c232
*+ bl_0_232 br_0_232 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c232
*+ bl_0_232 br_0_232 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c232
*+ bl_0_232 br_0_232 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c232
*+ bl_0_232 br_0_232 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c232
*+ bl_0_232 br_0_232 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c232
*+ bl_0_232 br_0_232 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c232
*+ bl_0_232 br_0_232 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c232
*+ bl_0_232 br_0_232 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c232
*+ bl_0_232 br_0_232 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c232
*+ bl_0_232 br_0_232 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c232
*+ bl_0_232 br_0_232 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c232
*+ bl_0_232 br_0_232 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c232
*+ bl_0_232 br_0_232 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c232
*+ bl_0_232 br_0_232 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c232
*+ bl_0_232 br_0_232 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c232
*+ bl_0_232 br_0_232 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c232
*+ bl_0_232 br_0_232 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c232
*+ bl_0_232 br_0_232 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c232
*+ bl_0_232 br_0_232 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c232
*+ bl_0_232 br_0_232 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c232
*+ bl_0_232 br_0_232 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c232
*+ bl_0_232 br_0_232 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c232
*+ bl_0_232 br_0_232 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c232
*+ bl_0_232 br_0_232 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c232
*+ bl_0_232 br_0_232 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c232
*+ bl_0_232 br_0_232 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c232
*+ bl_0_232 br_0_232 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c232
*+ bl_0_232 br_0_232 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c232
*+ bl_0_232 br_0_232 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c232
*+ bl_0_232 br_0_232 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c232
*+ bl_0_232 br_0_232 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c232
*+ bl_0_232 br_0_232 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c232
*+ bl_0_232 br_0_232 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c232
*+ bl_0_232 br_0_232 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c232
*+ bl_0_232 br_0_232 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c232
*+ bl_0_232 br_0_232 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c232
*+ bl_0_232 br_0_232 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c232
*+ bl_0_232 br_0_232 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c232
*+ bl_0_232 br_0_232 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c232
*+ bl_0_232 br_0_232 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c232
*+ bl_0_232 br_0_232 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c232
*+ bl_0_232 br_0_232 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c232
*+ bl_0_232 br_0_232 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c232
*+ bl_0_232 br_0_232 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c232
*+ bl_0_232 br_0_232 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c232
*+ bl_0_232 br_0_232 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c232
*+ bl_0_232 br_0_232 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c232
*+ bl_0_232 br_0_232 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c232
*+ bl_0_232 br_0_232 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c232
*+ bl_0_232 br_0_232 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c232
*+ bl_0_232 br_0_232 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c232
*+ bl_0_232 br_0_232 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c232
*+ bl_0_232 br_0_232 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c232
*+ bl_0_232 br_0_232 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c232
*+ bl_0_232 br_0_232 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c232
*+ bl_0_232 br_0_232 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c232
*+ bl_0_232 br_0_232 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c232
*+ bl_0_232 br_0_232 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c232
*+ bl_0_232 br_0_232 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c232
*+ bl_0_232 br_0_232 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c232
*+ bl_0_232 br_0_232 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c232
*+ bl_0_232 br_0_232 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c232
*+ bl_0_232 br_0_232 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c232
*+ bl_0_232 br_0_232 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c232
*+ bl_0_232 br_0_232 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c232
*+ bl_0_232 br_0_232 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c232
*+ bl_0_232 br_0_232 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c232
*+ bl_0_232 br_0_232 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c232
*+ bl_0_232 br_0_232 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c232
*+ bl_0_232 br_0_232 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c232
*+ bl_0_232 br_0_232 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c232
*+ bl_0_232 br_0_232 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c232
*+ bl_0_232 br_0_232 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c232
*+ bl_0_232 br_0_232 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c232
*+ bl_0_232 br_0_232 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c232
*+ bl_0_232 br_0_232 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c232
*+ bl_0_232 br_0_232 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c232
*+ bl_0_232 br_0_232 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c232
*+ bl_0_232 br_0_232 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c232
*+ bl_0_232 br_0_232 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c232
*+ bl_0_232 br_0_232 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c232
*+ bl_0_232 br_0_232 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c232
*+ bl_0_232 br_0_232 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c232
*+ bl_0_232 br_0_232 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c232
*+ bl_0_232 br_0_232 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c232
*+ bl_0_232 br_0_232 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c232
*+ bl_0_232 br_0_232 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c232
*+ bl_0_232 br_0_232 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c232
*+ bl_0_232 br_0_232 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c232
*+ bl_0_232 br_0_232 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c232
*+ bl_0_232 br_0_232 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c232
*+ bl_0_232 br_0_232 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c232
*+ bl_0_232 br_0_232 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c232
*+ bl_0_232 br_0_232 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c232
*+ bl_0_232 br_0_232 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c232
*+ bl_0_232 br_0_232 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c232
*+ bl_0_232 br_0_232 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c232
*+ bl_0_232 br_0_232 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c232
*+ bl_0_232 br_0_232 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c232
*+ bl_0_232 br_0_232 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c232
*+ bl_0_232 br_0_232 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c232
*+ bl_0_232 br_0_232 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c232
*+ bl_0_232 br_0_232 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c232
*+ bl_0_232 br_0_232 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c232
*+ bl_0_232 br_0_232 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c232
+ bl_0_232 br_0_232 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c233
+ bl_0_233 br_0_233 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c233
*+ bl_0_233 br_0_233 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c233
*+ bl_0_233 br_0_233 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c233
*+ bl_0_233 br_0_233 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c233
*+ bl_0_233 br_0_233 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c233
*+ bl_0_233 br_0_233 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c233
*+ bl_0_233 br_0_233 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c233
*+ bl_0_233 br_0_233 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c233
*+ bl_0_233 br_0_233 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c233
*+ bl_0_233 br_0_233 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c233
*+ bl_0_233 br_0_233 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c233
*+ bl_0_233 br_0_233 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c233
*+ bl_0_233 br_0_233 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c233
*+ bl_0_233 br_0_233 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c233
*+ bl_0_233 br_0_233 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c233
*+ bl_0_233 br_0_233 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c233
*+ bl_0_233 br_0_233 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c233
*+ bl_0_233 br_0_233 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c233
*+ bl_0_233 br_0_233 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c233
*+ bl_0_233 br_0_233 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c233
*+ bl_0_233 br_0_233 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c233
*+ bl_0_233 br_0_233 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c233
*+ bl_0_233 br_0_233 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c233
*+ bl_0_233 br_0_233 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c233
*+ bl_0_233 br_0_233 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c233
*+ bl_0_233 br_0_233 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c233
*+ bl_0_233 br_0_233 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c233
*+ bl_0_233 br_0_233 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c233
*+ bl_0_233 br_0_233 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c233
*+ bl_0_233 br_0_233 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c233
*+ bl_0_233 br_0_233 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c233
*+ bl_0_233 br_0_233 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c233
*+ bl_0_233 br_0_233 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c233
*+ bl_0_233 br_0_233 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c233
*+ bl_0_233 br_0_233 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c233
*+ bl_0_233 br_0_233 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c233
*+ bl_0_233 br_0_233 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c233
*+ bl_0_233 br_0_233 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c233
*+ bl_0_233 br_0_233 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c233
*+ bl_0_233 br_0_233 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c233
*+ bl_0_233 br_0_233 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c233
*+ bl_0_233 br_0_233 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c233
*+ bl_0_233 br_0_233 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c233
*+ bl_0_233 br_0_233 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c233
*+ bl_0_233 br_0_233 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c233
*+ bl_0_233 br_0_233 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c233
*+ bl_0_233 br_0_233 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c233
*+ bl_0_233 br_0_233 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c233
*+ bl_0_233 br_0_233 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c233
*+ bl_0_233 br_0_233 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c233
*+ bl_0_233 br_0_233 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c233
*+ bl_0_233 br_0_233 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c233
*+ bl_0_233 br_0_233 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c233
*+ bl_0_233 br_0_233 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c233
*+ bl_0_233 br_0_233 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c233
*+ bl_0_233 br_0_233 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c233
*+ bl_0_233 br_0_233 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c233
*+ bl_0_233 br_0_233 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c233
*+ bl_0_233 br_0_233 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c233
*+ bl_0_233 br_0_233 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c233
*+ bl_0_233 br_0_233 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c233
*+ bl_0_233 br_0_233 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c233
*+ bl_0_233 br_0_233 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c233
*+ bl_0_233 br_0_233 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c233
*+ bl_0_233 br_0_233 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c233
*+ bl_0_233 br_0_233 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c233
*+ bl_0_233 br_0_233 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c233
*+ bl_0_233 br_0_233 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c233
*+ bl_0_233 br_0_233 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c233
*+ bl_0_233 br_0_233 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c233
*+ bl_0_233 br_0_233 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c233
*+ bl_0_233 br_0_233 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c233
*+ bl_0_233 br_0_233 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c233
*+ bl_0_233 br_0_233 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c233
*+ bl_0_233 br_0_233 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c233
*+ bl_0_233 br_0_233 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c233
*+ bl_0_233 br_0_233 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c233
*+ bl_0_233 br_0_233 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c233
*+ bl_0_233 br_0_233 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c233
*+ bl_0_233 br_0_233 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c233
*+ bl_0_233 br_0_233 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c233
*+ bl_0_233 br_0_233 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c233
*+ bl_0_233 br_0_233 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c233
*+ bl_0_233 br_0_233 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c233
*+ bl_0_233 br_0_233 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c233
*+ bl_0_233 br_0_233 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c233
*+ bl_0_233 br_0_233 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c233
*+ bl_0_233 br_0_233 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c233
*+ bl_0_233 br_0_233 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c233
*+ bl_0_233 br_0_233 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c233
*+ bl_0_233 br_0_233 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c233
*+ bl_0_233 br_0_233 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c233
*+ bl_0_233 br_0_233 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c233
*+ bl_0_233 br_0_233 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c233
*+ bl_0_233 br_0_233 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c233
*+ bl_0_233 br_0_233 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c233
*+ bl_0_233 br_0_233 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c233
*+ bl_0_233 br_0_233 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c233
*+ bl_0_233 br_0_233 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c233
*+ bl_0_233 br_0_233 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c233
*+ bl_0_233 br_0_233 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c233
*+ bl_0_233 br_0_233 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c233
*+ bl_0_233 br_0_233 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c233
*+ bl_0_233 br_0_233 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c233
*+ bl_0_233 br_0_233 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c233
*+ bl_0_233 br_0_233 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c233
*+ bl_0_233 br_0_233 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c233
*+ bl_0_233 br_0_233 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c233
*+ bl_0_233 br_0_233 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c233
*+ bl_0_233 br_0_233 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c233
*+ bl_0_233 br_0_233 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c233
*+ bl_0_233 br_0_233 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c233
*+ bl_0_233 br_0_233 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c233
*+ bl_0_233 br_0_233 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c233
*+ bl_0_233 br_0_233 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c233
*+ bl_0_233 br_0_233 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c233
*+ bl_0_233 br_0_233 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c233
*+ bl_0_233 br_0_233 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c233
*+ bl_0_233 br_0_233 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c233
*+ bl_0_233 br_0_233 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c233
*+ bl_0_233 br_0_233 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c233
*+ bl_0_233 br_0_233 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c233
*+ bl_0_233 br_0_233 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c233
*+ bl_0_233 br_0_233 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c233
*+ bl_0_233 br_0_233 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c233
*+ bl_0_233 br_0_233 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c233
*+ bl_0_233 br_0_233 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c233
+ bl_0_233 br_0_233 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c234
+ bl_0_234 br_0_234 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c234
*+ bl_0_234 br_0_234 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c234
*+ bl_0_234 br_0_234 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c234
*+ bl_0_234 br_0_234 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c234
*+ bl_0_234 br_0_234 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c234
*+ bl_0_234 br_0_234 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c234
*+ bl_0_234 br_0_234 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c234
*+ bl_0_234 br_0_234 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c234
*+ bl_0_234 br_0_234 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c234
*+ bl_0_234 br_0_234 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c234
*+ bl_0_234 br_0_234 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c234
*+ bl_0_234 br_0_234 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c234
*+ bl_0_234 br_0_234 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c234
*+ bl_0_234 br_0_234 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c234
*+ bl_0_234 br_0_234 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c234
*+ bl_0_234 br_0_234 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c234
*+ bl_0_234 br_0_234 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c234
*+ bl_0_234 br_0_234 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c234
*+ bl_0_234 br_0_234 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c234
*+ bl_0_234 br_0_234 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c234
*+ bl_0_234 br_0_234 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c234
*+ bl_0_234 br_0_234 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c234
*+ bl_0_234 br_0_234 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c234
*+ bl_0_234 br_0_234 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c234
*+ bl_0_234 br_0_234 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c234
*+ bl_0_234 br_0_234 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c234
*+ bl_0_234 br_0_234 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c234
*+ bl_0_234 br_0_234 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c234
*+ bl_0_234 br_0_234 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c234
*+ bl_0_234 br_0_234 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c234
*+ bl_0_234 br_0_234 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c234
*+ bl_0_234 br_0_234 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c234
*+ bl_0_234 br_0_234 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c234
*+ bl_0_234 br_0_234 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c234
*+ bl_0_234 br_0_234 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c234
*+ bl_0_234 br_0_234 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c234
*+ bl_0_234 br_0_234 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c234
*+ bl_0_234 br_0_234 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c234
*+ bl_0_234 br_0_234 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c234
*+ bl_0_234 br_0_234 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c234
*+ bl_0_234 br_0_234 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c234
*+ bl_0_234 br_0_234 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c234
*+ bl_0_234 br_0_234 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c234
*+ bl_0_234 br_0_234 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c234
*+ bl_0_234 br_0_234 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c234
*+ bl_0_234 br_0_234 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c234
*+ bl_0_234 br_0_234 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c234
*+ bl_0_234 br_0_234 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c234
*+ bl_0_234 br_0_234 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c234
*+ bl_0_234 br_0_234 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c234
*+ bl_0_234 br_0_234 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c234
*+ bl_0_234 br_0_234 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c234
*+ bl_0_234 br_0_234 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c234
*+ bl_0_234 br_0_234 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c234
*+ bl_0_234 br_0_234 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c234
*+ bl_0_234 br_0_234 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c234
*+ bl_0_234 br_0_234 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c234
*+ bl_0_234 br_0_234 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c234
*+ bl_0_234 br_0_234 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c234
*+ bl_0_234 br_0_234 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c234
*+ bl_0_234 br_0_234 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c234
*+ bl_0_234 br_0_234 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c234
*+ bl_0_234 br_0_234 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c234
*+ bl_0_234 br_0_234 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c234
*+ bl_0_234 br_0_234 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c234
*+ bl_0_234 br_0_234 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c234
*+ bl_0_234 br_0_234 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c234
*+ bl_0_234 br_0_234 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c234
*+ bl_0_234 br_0_234 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c234
*+ bl_0_234 br_0_234 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c234
*+ bl_0_234 br_0_234 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c234
*+ bl_0_234 br_0_234 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c234
*+ bl_0_234 br_0_234 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c234
*+ bl_0_234 br_0_234 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c234
*+ bl_0_234 br_0_234 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c234
*+ bl_0_234 br_0_234 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c234
*+ bl_0_234 br_0_234 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c234
*+ bl_0_234 br_0_234 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c234
*+ bl_0_234 br_0_234 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c234
*+ bl_0_234 br_0_234 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c234
*+ bl_0_234 br_0_234 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c234
*+ bl_0_234 br_0_234 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c234
*+ bl_0_234 br_0_234 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c234
*+ bl_0_234 br_0_234 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c234
*+ bl_0_234 br_0_234 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c234
*+ bl_0_234 br_0_234 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c234
*+ bl_0_234 br_0_234 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c234
*+ bl_0_234 br_0_234 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c234
*+ bl_0_234 br_0_234 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c234
*+ bl_0_234 br_0_234 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c234
*+ bl_0_234 br_0_234 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c234
*+ bl_0_234 br_0_234 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c234
*+ bl_0_234 br_0_234 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c234
*+ bl_0_234 br_0_234 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c234
*+ bl_0_234 br_0_234 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c234
*+ bl_0_234 br_0_234 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c234
*+ bl_0_234 br_0_234 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c234
*+ bl_0_234 br_0_234 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c234
*+ bl_0_234 br_0_234 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c234
*+ bl_0_234 br_0_234 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c234
*+ bl_0_234 br_0_234 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c234
*+ bl_0_234 br_0_234 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c234
*+ bl_0_234 br_0_234 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c234
*+ bl_0_234 br_0_234 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c234
*+ bl_0_234 br_0_234 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c234
*+ bl_0_234 br_0_234 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c234
*+ bl_0_234 br_0_234 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c234
*+ bl_0_234 br_0_234 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c234
*+ bl_0_234 br_0_234 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c234
*+ bl_0_234 br_0_234 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c234
*+ bl_0_234 br_0_234 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c234
*+ bl_0_234 br_0_234 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c234
*+ bl_0_234 br_0_234 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c234
*+ bl_0_234 br_0_234 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c234
*+ bl_0_234 br_0_234 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c234
*+ bl_0_234 br_0_234 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c234
*+ bl_0_234 br_0_234 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c234
*+ bl_0_234 br_0_234 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c234
*+ bl_0_234 br_0_234 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c234
*+ bl_0_234 br_0_234 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c234
*+ bl_0_234 br_0_234 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c234
*+ bl_0_234 br_0_234 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c234
*+ bl_0_234 br_0_234 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c234
*+ bl_0_234 br_0_234 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c234
*+ bl_0_234 br_0_234 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c234
*+ bl_0_234 br_0_234 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c234
*+ bl_0_234 br_0_234 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c234
+ bl_0_234 br_0_234 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c235
+ bl_0_235 br_0_235 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c235
*+ bl_0_235 br_0_235 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c235
*+ bl_0_235 br_0_235 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c235
*+ bl_0_235 br_0_235 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c235
*+ bl_0_235 br_0_235 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c235
*+ bl_0_235 br_0_235 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c235
*+ bl_0_235 br_0_235 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c235
*+ bl_0_235 br_0_235 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c235
*+ bl_0_235 br_0_235 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c235
*+ bl_0_235 br_0_235 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c235
*+ bl_0_235 br_0_235 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c235
*+ bl_0_235 br_0_235 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c235
*+ bl_0_235 br_0_235 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c235
*+ bl_0_235 br_0_235 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c235
*+ bl_0_235 br_0_235 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c235
*+ bl_0_235 br_0_235 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c235
*+ bl_0_235 br_0_235 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c235
*+ bl_0_235 br_0_235 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c235
*+ bl_0_235 br_0_235 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c235
*+ bl_0_235 br_0_235 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c235
*+ bl_0_235 br_0_235 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c235
*+ bl_0_235 br_0_235 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c235
*+ bl_0_235 br_0_235 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c235
*+ bl_0_235 br_0_235 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c235
*+ bl_0_235 br_0_235 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c235
*+ bl_0_235 br_0_235 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c235
*+ bl_0_235 br_0_235 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c235
*+ bl_0_235 br_0_235 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c235
*+ bl_0_235 br_0_235 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c235
*+ bl_0_235 br_0_235 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c235
*+ bl_0_235 br_0_235 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c235
*+ bl_0_235 br_0_235 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c235
*+ bl_0_235 br_0_235 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c235
*+ bl_0_235 br_0_235 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c235
*+ bl_0_235 br_0_235 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c235
*+ bl_0_235 br_0_235 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c235
*+ bl_0_235 br_0_235 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c235
*+ bl_0_235 br_0_235 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c235
*+ bl_0_235 br_0_235 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c235
*+ bl_0_235 br_0_235 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c235
*+ bl_0_235 br_0_235 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c235
*+ bl_0_235 br_0_235 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c235
*+ bl_0_235 br_0_235 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c235
*+ bl_0_235 br_0_235 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c235
*+ bl_0_235 br_0_235 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c235
*+ bl_0_235 br_0_235 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c235
*+ bl_0_235 br_0_235 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c235
*+ bl_0_235 br_0_235 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c235
*+ bl_0_235 br_0_235 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c235
*+ bl_0_235 br_0_235 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c235
*+ bl_0_235 br_0_235 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c235
*+ bl_0_235 br_0_235 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c235
*+ bl_0_235 br_0_235 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c235
*+ bl_0_235 br_0_235 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c235
*+ bl_0_235 br_0_235 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c235
*+ bl_0_235 br_0_235 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c235
*+ bl_0_235 br_0_235 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c235
*+ bl_0_235 br_0_235 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c235
*+ bl_0_235 br_0_235 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c235
*+ bl_0_235 br_0_235 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c235
*+ bl_0_235 br_0_235 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c235
*+ bl_0_235 br_0_235 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c235
*+ bl_0_235 br_0_235 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c235
*+ bl_0_235 br_0_235 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c235
*+ bl_0_235 br_0_235 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c235
*+ bl_0_235 br_0_235 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c235
*+ bl_0_235 br_0_235 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c235
*+ bl_0_235 br_0_235 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c235
*+ bl_0_235 br_0_235 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c235
*+ bl_0_235 br_0_235 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c235
*+ bl_0_235 br_0_235 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c235
*+ bl_0_235 br_0_235 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c235
*+ bl_0_235 br_0_235 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c235
*+ bl_0_235 br_0_235 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c235
*+ bl_0_235 br_0_235 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c235
*+ bl_0_235 br_0_235 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c235
*+ bl_0_235 br_0_235 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c235
*+ bl_0_235 br_0_235 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c235
*+ bl_0_235 br_0_235 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c235
*+ bl_0_235 br_0_235 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c235
*+ bl_0_235 br_0_235 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c235
*+ bl_0_235 br_0_235 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c235
*+ bl_0_235 br_0_235 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c235
*+ bl_0_235 br_0_235 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c235
*+ bl_0_235 br_0_235 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c235
*+ bl_0_235 br_0_235 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c235
*+ bl_0_235 br_0_235 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c235
*+ bl_0_235 br_0_235 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c235
*+ bl_0_235 br_0_235 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c235
*+ bl_0_235 br_0_235 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c235
*+ bl_0_235 br_0_235 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c235
*+ bl_0_235 br_0_235 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c235
*+ bl_0_235 br_0_235 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c235
*+ bl_0_235 br_0_235 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c235
*+ bl_0_235 br_0_235 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c235
*+ bl_0_235 br_0_235 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c235
*+ bl_0_235 br_0_235 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c235
*+ bl_0_235 br_0_235 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c235
*+ bl_0_235 br_0_235 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c235
*+ bl_0_235 br_0_235 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c235
*+ bl_0_235 br_0_235 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c235
*+ bl_0_235 br_0_235 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c235
*+ bl_0_235 br_0_235 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c235
*+ bl_0_235 br_0_235 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c235
*+ bl_0_235 br_0_235 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c235
*+ bl_0_235 br_0_235 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c235
*+ bl_0_235 br_0_235 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c235
*+ bl_0_235 br_0_235 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c235
*+ bl_0_235 br_0_235 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c235
*+ bl_0_235 br_0_235 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c235
*+ bl_0_235 br_0_235 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c235
*+ bl_0_235 br_0_235 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c235
*+ bl_0_235 br_0_235 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c235
*+ bl_0_235 br_0_235 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c235
*+ bl_0_235 br_0_235 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c235
*+ bl_0_235 br_0_235 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c235
*+ bl_0_235 br_0_235 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c235
*+ bl_0_235 br_0_235 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c235
*+ bl_0_235 br_0_235 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c235
*+ bl_0_235 br_0_235 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c235
*+ bl_0_235 br_0_235 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c235
*+ bl_0_235 br_0_235 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c235
*+ bl_0_235 br_0_235 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c235
*+ bl_0_235 br_0_235 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c235
*+ bl_0_235 br_0_235 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c235
*+ bl_0_235 br_0_235 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c235
*+ bl_0_235 br_0_235 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c235
+ bl_0_235 br_0_235 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c236
+ bl_0_236 br_0_236 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c236
*+ bl_0_236 br_0_236 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c236
*+ bl_0_236 br_0_236 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c236
*+ bl_0_236 br_0_236 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c236
*+ bl_0_236 br_0_236 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c236
*+ bl_0_236 br_0_236 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c236
*+ bl_0_236 br_0_236 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c236
*+ bl_0_236 br_0_236 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c236
*+ bl_0_236 br_0_236 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c236
*+ bl_0_236 br_0_236 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c236
*+ bl_0_236 br_0_236 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c236
*+ bl_0_236 br_0_236 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c236
*+ bl_0_236 br_0_236 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c236
*+ bl_0_236 br_0_236 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c236
*+ bl_0_236 br_0_236 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c236
*+ bl_0_236 br_0_236 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c236
*+ bl_0_236 br_0_236 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c236
*+ bl_0_236 br_0_236 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c236
*+ bl_0_236 br_0_236 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c236
*+ bl_0_236 br_0_236 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c236
*+ bl_0_236 br_0_236 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c236
*+ bl_0_236 br_0_236 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c236
*+ bl_0_236 br_0_236 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c236
*+ bl_0_236 br_0_236 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c236
*+ bl_0_236 br_0_236 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c236
*+ bl_0_236 br_0_236 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c236
*+ bl_0_236 br_0_236 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c236
*+ bl_0_236 br_0_236 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c236
*+ bl_0_236 br_0_236 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c236
*+ bl_0_236 br_0_236 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c236
*+ bl_0_236 br_0_236 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c236
*+ bl_0_236 br_0_236 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c236
*+ bl_0_236 br_0_236 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c236
*+ bl_0_236 br_0_236 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c236
*+ bl_0_236 br_0_236 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c236
*+ bl_0_236 br_0_236 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c236
*+ bl_0_236 br_0_236 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c236
*+ bl_0_236 br_0_236 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c236
*+ bl_0_236 br_0_236 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c236
*+ bl_0_236 br_0_236 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c236
*+ bl_0_236 br_0_236 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c236
*+ bl_0_236 br_0_236 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c236
*+ bl_0_236 br_0_236 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c236
*+ bl_0_236 br_0_236 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c236
*+ bl_0_236 br_0_236 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c236
*+ bl_0_236 br_0_236 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c236
*+ bl_0_236 br_0_236 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c236
*+ bl_0_236 br_0_236 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c236
*+ bl_0_236 br_0_236 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c236
*+ bl_0_236 br_0_236 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c236
*+ bl_0_236 br_0_236 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c236
*+ bl_0_236 br_0_236 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c236
*+ bl_0_236 br_0_236 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c236
*+ bl_0_236 br_0_236 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c236
*+ bl_0_236 br_0_236 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c236
*+ bl_0_236 br_0_236 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c236
*+ bl_0_236 br_0_236 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c236
*+ bl_0_236 br_0_236 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c236
*+ bl_0_236 br_0_236 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c236
*+ bl_0_236 br_0_236 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c236
*+ bl_0_236 br_0_236 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c236
*+ bl_0_236 br_0_236 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c236
*+ bl_0_236 br_0_236 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c236
*+ bl_0_236 br_0_236 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c236
*+ bl_0_236 br_0_236 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c236
*+ bl_0_236 br_0_236 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c236
*+ bl_0_236 br_0_236 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c236
*+ bl_0_236 br_0_236 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c236
*+ bl_0_236 br_0_236 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c236
*+ bl_0_236 br_0_236 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c236
*+ bl_0_236 br_0_236 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c236
*+ bl_0_236 br_0_236 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c236
*+ bl_0_236 br_0_236 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c236
*+ bl_0_236 br_0_236 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c236
*+ bl_0_236 br_0_236 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c236
*+ bl_0_236 br_0_236 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c236
*+ bl_0_236 br_0_236 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c236
*+ bl_0_236 br_0_236 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c236
*+ bl_0_236 br_0_236 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c236
*+ bl_0_236 br_0_236 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c236
*+ bl_0_236 br_0_236 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c236
*+ bl_0_236 br_0_236 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c236
*+ bl_0_236 br_0_236 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c236
*+ bl_0_236 br_0_236 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c236
*+ bl_0_236 br_0_236 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c236
*+ bl_0_236 br_0_236 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c236
*+ bl_0_236 br_0_236 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c236
*+ bl_0_236 br_0_236 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c236
*+ bl_0_236 br_0_236 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c236
*+ bl_0_236 br_0_236 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c236
*+ bl_0_236 br_0_236 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c236
*+ bl_0_236 br_0_236 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c236
*+ bl_0_236 br_0_236 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c236
*+ bl_0_236 br_0_236 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c236
*+ bl_0_236 br_0_236 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c236
*+ bl_0_236 br_0_236 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c236
*+ bl_0_236 br_0_236 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c236
*+ bl_0_236 br_0_236 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c236
*+ bl_0_236 br_0_236 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c236
*+ bl_0_236 br_0_236 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c236
*+ bl_0_236 br_0_236 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c236
*+ bl_0_236 br_0_236 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c236
*+ bl_0_236 br_0_236 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c236
*+ bl_0_236 br_0_236 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c236
*+ bl_0_236 br_0_236 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c236
*+ bl_0_236 br_0_236 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c236
*+ bl_0_236 br_0_236 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c236
*+ bl_0_236 br_0_236 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c236
*+ bl_0_236 br_0_236 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c236
*+ bl_0_236 br_0_236 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c236
*+ bl_0_236 br_0_236 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c236
*+ bl_0_236 br_0_236 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c236
*+ bl_0_236 br_0_236 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c236
*+ bl_0_236 br_0_236 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c236
*+ bl_0_236 br_0_236 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c236
*+ bl_0_236 br_0_236 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c236
*+ bl_0_236 br_0_236 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c236
*+ bl_0_236 br_0_236 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c236
*+ bl_0_236 br_0_236 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c236
*+ bl_0_236 br_0_236 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c236
*+ bl_0_236 br_0_236 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c236
*+ bl_0_236 br_0_236 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c236
*+ bl_0_236 br_0_236 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c236
*+ bl_0_236 br_0_236 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c236
*+ bl_0_236 br_0_236 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c236
*+ bl_0_236 br_0_236 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c236
*+ bl_0_236 br_0_236 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c236
+ bl_0_236 br_0_236 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c237
+ bl_0_237 br_0_237 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c237
*+ bl_0_237 br_0_237 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c237
*+ bl_0_237 br_0_237 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c237
*+ bl_0_237 br_0_237 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c237
*+ bl_0_237 br_0_237 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c237
*+ bl_0_237 br_0_237 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c237
*+ bl_0_237 br_0_237 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c237
*+ bl_0_237 br_0_237 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c237
*+ bl_0_237 br_0_237 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c237
*+ bl_0_237 br_0_237 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c237
*+ bl_0_237 br_0_237 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c237
*+ bl_0_237 br_0_237 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c237
*+ bl_0_237 br_0_237 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c237
*+ bl_0_237 br_0_237 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c237
*+ bl_0_237 br_0_237 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c237
*+ bl_0_237 br_0_237 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c237
*+ bl_0_237 br_0_237 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c237
*+ bl_0_237 br_0_237 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c237
*+ bl_0_237 br_0_237 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c237
*+ bl_0_237 br_0_237 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c237
*+ bl_0_237 br_0_237 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c237
*+ bl_0_237 br_0_237 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c237
*+ bl_0_237 br_0_237 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c237
*+ bl_0_237 br_0_237 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c237
*+ bl_0_237 br_0_237 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c237
*+ bl_0_237 br_0_237 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c237
*+ bl_0_237 br_0_237 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c237
*+ bl_0_237 br_0_237 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c237
*+ bl_0_237 br_0_237 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c237
*+ bl_0_237 br_0_237 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c237
*+ bl_0_237 br_0_237 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c237
*+ bl_0_237 br_0_237 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c237
*+ bl_0_237 br_0_237 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c237
*+ bl_0_237 br_0_237 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c237
*+ bl_0_237 br_0_237 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c237
*+ bl_0_237 br_0_237 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c237
*+ bl_0_237 br_0_237 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c237
*+ bl_0_237 br_0_237 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c237
*+ bl_0_237 br_0_237 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c237
*+ bl_0_237 br_0_237 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c237
*+ bl_0_237 br_0_237 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c237
*+ bl_0_237 br_0_237 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c237
*+ bl_0_237 br_0_237 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c237
*+ bl_0_237 br_0_237 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c237
*+ bl_0_237 br_0_237 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c237
*+ bl_0_237 br_0_237 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c237
*+ bl_0_237 br_0_237 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c237
*+ bl_0_237 br_0_237 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c237
*+ bl_0_237 br_0_237 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c237
*+ bl_0_237 br_0_237 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c237
*+ bl_0_237 br_0_237 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c237
*+ bl_0_237 br_0_237 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c237
*+ bl_0_237 br_0_237 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c237
*+ bl_0_237 br_0_237 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c237
*+ bl_0_237 br_0_237 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c237
*+ bl_0_237 br_0_237 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c237
*+ bl_0_237 br_0_237 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c237
*+ bl_0_237 br_0_237 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c237
*+ bl_0_237 br_0_237 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c237
*+ bl_0_237 br_0_237 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c237
*+ bl_0_237 br_0_237 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c237
*+ bl_0_237 br_0_237 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c237
*+ bl_0_237 br_0_237 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c237
*+ bl_0_237 br_0_237 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c237
*+ bl_0_237 br_0_237 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c237
*+ bl_0_237 br_0_237 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c237
*+ bl_0_237 br_0_237 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c237
*+ bl_0_237 br_0_237 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c237
*+ bl_0_237 br_0_237 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c237
*+ bl_0_237 br_0_237 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c237
*+ bl_0_237 br_0_237 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c237
*+ bl_0_237 br_0_237 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c237
*+ bl_0_237 br_0_237 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c237
*+ bl_0_237 br_0_237 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c237
*+ bl_0_237 br_0_237 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c237
*+ bl_0_237 br_0_237 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c237
*+ bl_0_237 br_0_237 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c237
*+ bl_0_237 br_0_237 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c237
*+ bl_0_237 br_0_237 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c237
*+ bl_0_237 br_0_237 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c237
*+ bl_0_237 br_0_237 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c237
*+ bl_0_237 br_0_237 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c237
*+ bl_0_237 br_0_237 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c237
*+ bl_0_237 br_0_237 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c237
*+ bl_0_237 br_0_237 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c237
*+ bl_0_237 br_0_237 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c237
*+ bl_0_237 br_0_237 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c237
*+ bl_0_237 br_0_237 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c237
*+ bl_0_237 br_0_237 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c237
*+ bl_0_237 br_0_237 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c237
*+ bl_0_237 br_0_237 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c237
*+ bl_0_237 br_0_237 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c237
*+ bl_0_237 br_0_237 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c237
*+ bl_0_237 br_0_237 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c237
*+ bl_0_237 br_0_237 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c237
*+ bl_0_237 br_0_237 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c237
*+ bl_0_237 br_0_237 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c237
*+ bl_0_237 br_0_237 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c237
*+ bl_0_237 br_0_237 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c237
*+ bl_0_237 br_0_237 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c237
*+ bl_0_237 br_0_237 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c237
*+ bl_0_237 br_0_237 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c237
*+ bl_0_237 br_0_237 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c237
*+ bl_0_237 br_0_237 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c237
*+ bl_0_237 br_0_237 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c237
*+ bl_0_237 br_0_237 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c237
*+ bl_0_237 br_0_237 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c237
*+ bl_0_237 br_0_237 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c237
*+ bl_0_237 br_0_237 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c237
*+ bl_0_237 br_0_237 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c237
*+ bl_0_237 br_0_237 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c237
*+ bl_0_237 br_0_237 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c237
*+ bl_0_237 br_0_237 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c237
*+ bl_0_237 br_0_237 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c237
*+ bl_0_237 br_0_237 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c237
*+ bl_0_237 br_0_237 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c237
*+ bl_0_237 br_0_237 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c237
*+ bl_0_237 br_0_237 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c237
*+ bl_0_237 br_0_237 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c237
*+ bl_0_237 br_0_237 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c237
*+ bl_0_237 br_0_237 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c237
*+ bl_0_237 br_0_237 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c237
*+ bl_0_237 br_0_237 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c237
*+ bl_0_237 br_0_237 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c237
*+ bl_0_237 br_0_237 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c237
*+ bl_0_237 br_0_237 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c237
*+ bl_0_237 br_0_237 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c237
+ bl_0_237 br_0_237 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c238
+ bl_0_238 br_0_238 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c238
*+ bl_0_238 br_0_238 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c238
*+ bl_0_238 br_0_238 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c238
*+ bl_0_238 br_0_238 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c238
*+ bl_0_238 br_0_238 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c238
*+ bl_0_238 br_0_238 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c238
*+ bl_0_238 br_0_238 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c238
*+ bl_0_238 br_0_238 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c238
*+ bl_0_238 br_0_238 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c238
*+ bl_0_238 br_0_238 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c238
*+ bl_0_238 br_0_238 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c238
*+ bl_0_238 br_0_238 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c238
*+ bl_0_238 br_0_238 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c238
*+ bl_0_238 br_0_238 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c238
*+ bl_0_238 br_0_238 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c238
*+ bl_0_238 br_0_238 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c238
*+ bl_0_238 br_0_238 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c238
*+ bl_0_238 br_0_238 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c238
*+ bl_0_238 br_0_238 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c238
*+ bl_0_238 br_0_238 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c238
*+ bl_0_238 br_0_238 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c238
*+ bl_0_238 br_0_238 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c238
*+ bl_0_238 br_0_238 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c238
*+ bl_0_238 br_0_238 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c238
*+ bl_0_238 br_0_238 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c238
*+ bl_0_238 br_0_238 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c238
*+ bl_0_238 br_0_238 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c238
*+ bl_0_238 br_0_238 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c238
*+ bl_0_238 br_0_238 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c238
*+ bl_0_238 br_0_238 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c238
*+ bl_0_238 br_0_238 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c238
*+ bl_0_238 br_0_238 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c238
*+ bl_0_238 br_0_238 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c238
*+ bl_0_238 br_0_238 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c238
*+ bl_0_238 br_0_238 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c238
*+ bl_0_238 br_0_238 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c238
*+ bl_0_238 br_0_238 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c238
*+ bl_0_238 br_0_238 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c238
*+ bl_0_238 br_0_238 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c238
*+ bl_0_238 br_0_238 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c238
*+ bl_0_238 br_0_238 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c238
*+ bl_0_238 br_0_238 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c238
*+ bl_0_238 br_0_238 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c238
*+ bl_0_238 br_0_238 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c238
*+ bl_0_238 br_0_238 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c238
*+ bl_0_238 br_0_238 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c238
*+ bl_0_238 br_0_238 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c238
*+ bl_0_238 br_0_238 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c238
*+ bl_0_238 br_0_238 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c238
*+ bl_0_238 br_0_238 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c238
*+ bl_0_238 br_0_238 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c238
*+ bl_0_238 br_0_238 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c238
*+ bl_0_238 br_0_238 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c238
*+ bl_0_238 br_0_238 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c238
*+ bl_0_238 br_0_238 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c238
*+ bl_0_238 br_0_238 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c238
*+ bl_0_238 br_0_238 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c238
*+ bl_0_238 br_0_238 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c238
*+ bl_0_238 br_0_238 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c238
*+ bl_0_238 br_0_238 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c238
*+ bl_0_238 br_0_238 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c238
*+ bl_0_238 br_0_238 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c238
*+ bl_0_238 br_0_238 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c238
*+ bl_0_238 br_0_238 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c238
*+ bl_0_238 br_0_238 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c238
*+ bl_0_238 br_0_238 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c238
*+ bl_0_238 br_0_238 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c238
*+ bl_0_238 br_0_238 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c238
*+ bl_0_238 br_0_238 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c238
*+ bl_0_238 br_0_238 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c238
*+ bl_0_238 br_0_238 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c238
*+ bl_0_238 br_0_238 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c238
*+ bl_0_238 br_0_238 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c238
*+ bl_0_238 br_0_238 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c238
*+ bl_0_238 br_0_238 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c238
*+ bl_0_238 br_0_238 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c238
*+ bl_0_238 br_0_238 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c238
*+ bl_0_238 br_0_238 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c238
*+ bl_0_238 br_0_238 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c238
*+ bl_0_238 br_0_238 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c238
*+ bl_0_238 br_0_238 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c238
*+ bl_0_238 br_0_238 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c238
*+ bl_0_238 br_0_238 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c238
*+ bl_0_238 br_0_238 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c238
*+ bl_0_238 br_0_238 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c238
*+ bl_0_238 br_0_238 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c238
*+ bl_0_238 br_0_238 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c238
*+ bl_0_238 br_0_238 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c238
*+ bl_0_238 br_0_238 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c238
*+ bl_0_238 br_0_238 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c238
*+ bl_0_238 br_0_238 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c238
*+ bl_0_238 br_0_238 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c238
*+ bl_0_238 br_0_238 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c238
*+ bl_0_238 br_0_238 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c238
*+ bl_0_238 br_0_238 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c238
*+ bl_0_238 br_0_238 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c238
*+ bl_0_238 br_0_238 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c238
*+ bl_0_238 br_0_238 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c238
*+ bl_0_238 br_0_238 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c238
*+ bl_0_238 br_0_238 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c238
*+ bl_0_238 br_0_238 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c238
*+ bl_0_238 br_0_238 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c238
*+ bl_0_238 br_0_238 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c238
*+ bl_0_238 br_0_238 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c238
*+ bl_0_238 br_0_238 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c238
*+ bl_0_238 br_0_238 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c238
*+ bl_0_238 br_0_238 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c238
*+ bl_0_238 br_0_238 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c238
*+ bl_0_238 br_0_238 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c238
*+ bl_0_238 br_0_238 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c238
*+ bl_0_238 br_0_238 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c238
*+ bl_0_238 br_0_238 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c238
*+ bl_0_238 br_0_238 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c238
*+ bl_0_238 br_0_238 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c238
*+ bl_0_238 br_0_238 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c238
*+ bl_0_238 br_0_238 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c238
*+ bl_0_238 br_0_238 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c238
*+ bl_0_238 br_0_238 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c238
*+ bl_0_238 br_0_238 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c238
*+ bl_0_238 br_0_238 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c238
*+ bl_0_238 br_0_238 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c238
*+ bl_0_238 br_0_238 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c238
*+ bl_0_238 br_0_238 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c238
*+ bl_0_238 br_0_238 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c238
*+ bl_0_238 br_0_238 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c238
*+ bl_0_238 br_0_238 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c238
*+ bl_0_238 br_0_238 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c238
+ bl_0_238 br_0_238 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c239
+ bl_0_239 br_0_239 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c239
*+ bl_0_239 br_0_239 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c239
*+ bl_0_239 br_0_239 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c239
*+ bl_0_239 br_0_239 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c239
*+ bl_0_239 br_0_239 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c239
*+ bl_0_239 br_0_239 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c239
*+ bl_0_239 br_0_239 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c239
*+ bl_0_239 br_0_239 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c239
*+ bl_0_239 br_0_239 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c239
*+ bl_0_239 br_0_239 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c239
*+ bl_0_239 br_0_239 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c239
*+ bl_0_239 br_0_239 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c239
*+ bl_0_239 br_0_239 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c239
*+ bl_0_239 br_0_239 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c239
*+ bl_0_239 br_0_239 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c239
*+ bl_0_239 br_0_239 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c239
*+ bl_0_239 br_0_239 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c239
*+ bl_0_239 br_0_239 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c239
*+ bl_0_239 br_0_239 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c239
*+ bl_0_239 br_0_239 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c239
*+ bl_0_239 br_0_239 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c239
*+ bl_0_239 br_0_239 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c239
*+ bl_0_239 br_0_239 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c239
*+ bl_0_239 br_0_239 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c239
*+ bl_0_239 br_0_239 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c239
*+ bl_0_239 br_0_239 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c239
*+ bl_0_239 br_0_239 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c239
*+ bl_0_239 br_0_239 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c239
*+ bl_0_239 br_0_239 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c239
*+ bl_0_239 br_0_239 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c239
*+ bl_0_239 br_0_239 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c239
*+ bl_0_239 br_0_239 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c239
*+ bl_0_239 br_0_239 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c239
*+ bl_0_239 br_0_239 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c239
*+ bl_0_239 br_0_239 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c239
*+ bl_0_239 br_0_239 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c239
*+ bl_0_239 br_0_239 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c239
*+ bl_0_239 br_0_239 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c239
*+ bl_0_239 br_0_239 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c239
*+ bl_0_239 br_0_239 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c239
*+ bl_0_239 br_0_239 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c239
*+ bl_0_239 br_0_239 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c239
*+ bl_0_239 br_0_239 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c239
*+ bl_0_239 br_0_239 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c239
*+ bl_0_239 br_0_239 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c239
*+ bl_0_239 br_0_239 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c239
*+ bl_0_239 br_0_239 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c239
*+ bl_0_239 br_0_239 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c239
*+ bl_0_239 br_0_239 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c239
*+ bl_0_239 br_0_239 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c239
*+ bl_0_239 br_0_239 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c239
*+ bl_0_239 br_0_239 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c239
*+ bl_0_239 br_0_239 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c239
*+ bl_0_239 br_0_239 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c239
*+ bl_0_239 br_0_239 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c239
*+ bl_0_239 br_0_239 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c239
*+ bl_0_239 br_0_239 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c239
*+ bl_0_239 br_0_239 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c239
*+ bl_0_239 br_0_239 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c239
*+ bl_0_239 br_0_239 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c239
*+ bl_0_239 br_0_239 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c239
*+ bl_0_239 br_0_239 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c239
*+ bl_0_239 br_0_239 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c239
*+ bl_0_239 br_0_239 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c239
*+ bl_0_239 br_0_239 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c239
*+ bl_0_239 br_0_239 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c239
*+ bl_0_239 br_0_239 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c239
*+ bl_0_239 br_0_239 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c239
*+ bl_0_239 br_0_239 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c239
*+ bl_0_239 br_0_239 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c239
*+ bl_0_239 br_0_239 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c239
*+ bl_0_239 br_0_239 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c239
*+ bl_0_239 br_0_239 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c239
*+ bl_0_239 br_0_239 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c239
*+ bl_0_239 br_0_239 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c239
*+ bl_0_239 br_0_239 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c239
*+ bl_0_239 br_0_239 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c239
*+ bl_0_239 br_0_239 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c239
*+ bl_0_239 br_0_239 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c239
*+ bl_0_239 br_0_239 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c239
*+ bl_0_239 br_0_239 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c239
*+ bl_0_239 br_0_239 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c239
*+ bl_0_239 br_0_239 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c239
*+ bl_0_239 br_0_239 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c239
*+ bl_0_239 br_0_239 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c239
*+ bl_0_239 br_0_239 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c239
*+ bl_0_239 br_0_239 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c239
*+ bl_0_239 br_0_239 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c239
*+ bl_0_239 br_0_239 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c239
*+ bl_0_239 br_0_239 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c239
*+ bl_0_239 br_0_239 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c239
*+ bl_0_239 br_0_239 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c239
*+ bl_0_239 br_0_239 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c239
*+ bl_0_239 br_0_239 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c239
*+ bl_0_239 br_0_239 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c239
*+ bl_0_239 br_0_239 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c239
*+ bl_0_239 br_0_239 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c239
*+ bl_0_239 br_0_239 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c239
*+ bl_0_239 br_0_239 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c239
*+ bl_0_239 br_0_239 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c239
*+ bl_0_239 br_0_239 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c239
*+ bl_0_239 br_0_239 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c239
*+ bl_0_239 br_0_239 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c239
*+ bl_0_239 br_0_239 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c239
*+ bl_0_239 br_0_239 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c239
*+ bl_0_239 br_0_239 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c239
*+ bl_0_239 br_0_239 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c239
*+ bl_0_239 br_0_239 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c239
*+ bl_0_239 br_0_239 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c239
*+ bl_0_239 br_0_239 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c239
*+ bl_0_239 br_0_239 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c239
*+ bl_0_239 br_0_239 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c239
*+ bl_0_239 br_0_239 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c239
*+ bl_0_239 br_0_239 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c239
*+ bl_0_239 br_0_239 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c239
*+ bl_0_239 br_0_239 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c239
*+ bl_0_239 br_0_239 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c239
*+ bl_0_239 br_0_239 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c239
*+ bl_0_239 br_0_239 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c239
*+ bl_0_239 br_0_239 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c239
*+ bl_0_239 br_0_239 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c239
*+ bl_0_239 br_0_239 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c239
*+ bl_0_239 br_0_239 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c239
*+ bl_0_239 br_0_239 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c239
*+ bl_0_239 br_0_239 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c239
*+ bl_0_239 br_0_239 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c239
*+ bl_0_239 br_0_239 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c239
+ bl_0_239 br_0_239 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c240
+ bl_0_240 br_0_240 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c240
*+ bl_0_240 br_0_240 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c240
*+ bl_0_240 br_0_240 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c240
*+ bl_0_240 br_0_240 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c240
*+ bl_0_240 br_0_240 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c240
*+ bl_0_240 br_0_240 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c240
*+ bl_0_240 br_0_240 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c240
*+ bl_0_240 br_0_240 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c240
*+ bl_0_240 br_0_240 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c240
*+ bl_0_240 br_0_240 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c240
*+ bl_0_240 br_0_240 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c240
*+ bl_0_240 br_0_240 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c240
*+ bl_0_240 br_0_240 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c240
*+ bl_0_240 br_0_240 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c240
*+ bl_0_240 br_0_240 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c240
*+ bl_0_240 br_0_240 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c240
*+ bl_0_240 br_0_240 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c240
*+ bl_0_240 br_0_240 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c240
*+ bl_0_240 br_0_240 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c240
*+ bl_0_240 br_0_240 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c240
*+ bl_0_240 br_0_240 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c240
*+ bl_0_240 br_0_240 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c240
*+ bl_0_240 br_0_240 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c240
*+ bl_0_240 br_0_240 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c240
*+ bl_0_240 br_0_240 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c240
*+ bl_0_240 br_0_240 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c240
*+ bl_0_240 br_0_240 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c240
*+ bl_0_240 br_0_240 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c240
*+ bl_0_240 br_0_240 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c240
*+ bl_0_240 br_0_240 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c240
*+ bl_0_240 br_0_240 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c240
*+ bl_0_240 br_0_240 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c240
*+ bl_0_240 br_0_240 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c240
*+ bl_0_240 br_0_240 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c240
*+ bl_0_240 br_0_240 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c240
*+ bl_0_240 br_0_240 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c240
*+ bl_0_240 br_0_240 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c240
*+ bl_0_240 br_0_240 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c240
*+ bl_0_240 br_0_240 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c240
*+ bl_0_240 br_0_240 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c240
*+ bl_0_240 br_0_240 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c240
*+ bl_0_240 br_0_240 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c240
*+ bl_0_240 br_0_240 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c240
*+ bl_0_240 br_0_240 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c240
*+ bl_0_240 br_0_240 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c240
*+ bl_0_240 br_0_240 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c240
*+ bl_0_240 br_0_240 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c240
*+ bl_0_240 br_0_240 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c240
*+ bl_0_240 br_0_240 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c240
*+ bl_0_240 br_0_240 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c240
*+ bl_0_240 br_0_240 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c240
*+ bl_0_240 br_0_240 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c240
*+ bl_0_240 br_0_240 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c240
*+ bl_0_240 br_0_240 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c240
*+ bl_0_240 br_0_240 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c240
*+ bl_0_240 br_0_240 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c240
*+ bl_0_240 br_0_240 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c240
*+ bl_0_240 br_0_240 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c240
*+ bl_0_240 br_0_240 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c240
*+ bl_0_240 br_0_240 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c240
*+ bl_0_240 br_0_240 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c240
*+ bl_0_240 br_0_240 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c240
*+ bl_0_240 br_0_240 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c240
*+ bl_0_240 br_0_240 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c240
*+ bl_0_240 br_0_240 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c240
*+ bl_0_240 br_0_240 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c240
*+ bl_0_240 br_0_240 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c240
*+ bl_0_240 br_0_240 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c240
*+ bl_0_240 br_0_240 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c240
*+ bl_0_240 br_0_240 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c240
*+ bl_0_240 br_0_240 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c240
*+ bl_0_240 br_0_240 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c240
*+ bl_0_240 br_0_240 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c240
*+ bl_0_240 br_0_240 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c240
*+ bl_0_240 br_0_240 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c240
*+ bl_0_240 br_0_240 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c240
*+ bl_0_240 br_0_240 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c240
*+ bl_0_240 br_0_240 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c240
*+ bl_0_240 br_0_240 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c240
*+ bl_0_240 br_0_240 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c240
*+ bl_0_240 br_0_240 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c240
*+ bl_0_240 br_0_240 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c240
*+ bl_0_240 br_0_240 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c240
*+ bl_0_240 br_0_240 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c240
*+ bl_0_240 br_0_240 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c240
*+ bl_0_240 br_0_240 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c240
*+ bl_0_240 br_0_240 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c240
*+ bl_0_240 br_0_240 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c240
*+ bl_0_240 br_0_240 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c240
*+ bl_0_240 br_0_240 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c240
*+ bl_0_240 br_0_240 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c240
*+ bl_0_240 br_0_240 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c240
*+ bl_0_240 br_0_240 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c240
*+ bl_0_240 br_0_240 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c240
*+ bl_0_240 br_0_240 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c240
*+ bl_0_240 br_0_240 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c240
*+ bl_0_240 br_0_240 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c240
*+ bl_0_240 br_0_240 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c240
*+ bl_0_240 br_0_240 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c240
*+ bl_0_240 br_0_240 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c240
*+ bl_0_240 br_0_240 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c240
*+ bl_0_240 br_0_240 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c240
*+ bl_0_240 br_0_240 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c240
*+ bl_0_240 br_0_240 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c240
*+ bl_0_240 br_0_240 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c240
*+ bl_0_240 br_0_240 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c240
*+ bl_0_240 br_0_240 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c240
*+ bl_0_240 br_0_240 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c240
*+ bl_0_240 br_0_240 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c240
*+ bl_0_240 br_0_240 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c240
*+ bl_0_240 br_0_240 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c240
*+ bl_0_240 br_0_240 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c240
*+ bl_0_240 br_0_240 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c240
*+ bl_0_240 br_0_240 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c240
*+ bl_0_240 br_0_240 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c240
*+ bl_0_240 br_0_240 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c240
*+ bl_0_240 br_0_240 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c240
*+ bl_0_240 br_0_240 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c240
*+ bl_0_240 br_0_240 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c240
*+ bl_0_240 br_0_240 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c240
*+ bl_0_240 br_0_240 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c240
*+ bl_0_240 br_0_240 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c240
*+ bl_0_240 br_0_240 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c240
*+ bl_0_240 br_0_240 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c240
*+ bl_0_240 br_0_240 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c240
*+ bl_0_240 br_0_240 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c240
*+ bl_0_240 br_0_240 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c240
+ bl_0_240 br_0_240 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c241
+ bl_0_241 br_0_241 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c241
*+ bl_0_241 br_0_241 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c241
*+ bl_0_241 br_0_241 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c241
*+ bl_0_241 br_0_241 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c241
*+ bl_0_241 br_0_241 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c241
*+ bl_0_241 br_0_241 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c241
*+ bl_0_241 br_0_241 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c241
*+ bl_0_241 br_0_241 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c241
*+ bl_0_241 br_0_241 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c241
*+ bl_0_241 br_0_241 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c241
*+ bl_0_241 br_0_241 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c241
*+ bl_0_241 br_0_241 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c241
*+ bl_0_241 br_0_241 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c241
*+ bl_0_241 br_0_241 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c241
*+ bl_0_241 br_0_241 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c241
*+ bl_0_241 br_0_241 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c241
*+ bl_0_241 br_0_241 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c241
*+ bl_0_241 br_0_241 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c241
*+ bl_0_241 br_0_241 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c241
*+ bl_0_241 br_0_241 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c241
*+ bl_0_241 br_0_241 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c241
*+ bl_0_241 br_0_241 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c241
*+ bl_0_241 br_0_241 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c241
*+ bl_0_241 br_0_241 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c241
*+ bl_0_241 br_0_241 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c241
*+ bl_0_241 br_0_241 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c241
*+ bl_0_241 br_0_241 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c241
*+ bl_0_241 br_0_241 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c241
*+ bl_0_241 br_0_241 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c241
*+ bl_0_241 br_0_241 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c241
*+ bl_0_241 br_0_241 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c241
*+ bl_0_241 br_0_241 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c241
*+ bl_0_241 br_0_241 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c241
*+ bl_0_241 br_0_241 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c241
*+ bl_0_241 br_0_241 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c241
*+ bl_0_241 br_0_241 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c241
*+ bl_0_241 br_0_241 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c241
*+ bl_0_241 br_0_241 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c241
*+ bl_0_241 br_0_241 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c241
*+ bl_0_241 br_0_241 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c241
*+ bl_0_241 br_0_241 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c241
*+ bl_0_241 br_0_241 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c241
*+ bl_0_241 br_0_241 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c241
*+ bl_0_241 br_0_241 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c241
*+ bl_0_241 br_0_241 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c241
*+ bl_0_241 br_0_241 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c241
*+ bl_0_241 br_0_241 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c241
*+ bl_0_241 br_0_241 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c241
*+ bl_0_241 br_0_241 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c241
*+ bl_0_241 br_0_241 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c241
*+ bl_0_241 br_0_241 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c241
*+ bl_0_241 br_0_241 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c241
*+ bl_0_241 br_0_241 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c241
*+ bl_0_241 br_0_241 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c241
*+ bl_0_241 br_0_241 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c241
*+ bl_0_241 br_0_241 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c241
*+ bl_0_241 br_0_241 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c241
*+ bl_0_241 br_0_241 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c241
*+ bl_0_241 br_0_241 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c241
*+ bl_0_241 br_0_241 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c241
*+ bl_0_241 br_0_241 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c241
*+ bl_0_241 br_0_241 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c241
*+ bl_0_241 br_0_241 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c241
*+ bl_0_241 br_0_241 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c241
*+ bl_0_241 br_0_241 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c241
*+ bl_0_241 br_0_241 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c241
*+ bl_0_241 br_0_241 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c241
*+ bl_0_241 br_0_241 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c241
*+ bl_0_241 br_0_241 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c241
*+ bl_0_241 br_0_241 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c241
*+ bl_0_241 br_0_241 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c241
*+ bl_0_241 br_0_241 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c241
*+ bl_0_241 br_0_241 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c241
*+ bl_0_241 br_0_241 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c241
*+ bl_0_241 br_0_241 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c241
*+ bl_0_241 br_0_241 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c241
*+ bl_0_241 br_0_241 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c241
*+ bl_0_241 br_0_241 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c241
*+ bl_0_241 br_0_241 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c241
*+ bl_0_241 br_0_241 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c241
*+ bl_0_241 br_0_241 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c241
*+ bl_0_241 br_0_241 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c241
*+ bl_0_241 br_0_241 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c241
*+ bl_0_241 br_0_241 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c241
*+ bl_0_241 br_0_241 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c241
*+ bl_0_241 br_0_241 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c241
*+ bl_0_241 br_0_241 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c241
*+ bl_0_241 br_0_241 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c241
*+ bl_0_241 br_0_241 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c241
*+ bl_0_241 br_0_241 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c241
*+ bl_0_241 br_0_241 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c241
*+ bl_0_241 br_0_241 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c241
*+ bl_0_241 br_0_241 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c241
*+ bl_0_241 br_0_241 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c241
*+ bl_0_241 br_0_241 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c241
*+ bl_0_241 br_0_241 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c241
*+ bl_0_241 br_0_241 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c241
*+ bl_0_241 br_0_241 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c241
*+ bl_0_241 br_0_241 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c241
*+ bl_0_241 br_0_241 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c241
*+ bl_0_241 br_0_241 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c241
*+ bl_0_241 br_0_241 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c241
*+ bl_0_241 br_0_241 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c241
*+ bl_0_241 br_0_241 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c241
*+ bl_0_241 br_0_241 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c241
*+ bl_0_241 br_0_241 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c241
*+ bl_0_241 br_0_241 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c241
*+ bl_0_241 br_0_241 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c241
*+ bl_0_241 br_0_241 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c241
*+ bl_0_241 br_0_241 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c241
*+ bl_0_241 br_0_241 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c241
*+ bl_0_241 br_0_241 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c241
*+ bl_0_241 br_0_241 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c241
*+ bl_0_241 br_0_241 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c241
*+ bl_0_241 br_0_241 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c241
*+ bl_0_241 br_0_241 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c241
*+ bl_0_241 br_0_241 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c241
*+ bl_0_241 br_0_241 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c241
*+ bl_0_241 br_0_241 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c241
*+ bl_0_241 br_0_241 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c241
*+ bl_0_241 br_0_241 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c241
*+ bl_0_241 br_0_241 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c241
*+ bl_0_241 br_0_241 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c241
*+ bl_0_241 br_0_241 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c241
*+ bl_0_241 br_0_241 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c241
*+ bl_0_241 br_0_241 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c241
*+ bl_0_241 br_0_241 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c241
+ bl_0_241 br_0_241 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c242
+ bl_0_242 br_0_242 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c242
*+ bl_0_242 br_0_242 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c242
*+ bl_0_242 br_0_242 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c242
*+ bl_0_242 br_0_242 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c242
*+ bl_0_242 br_0_242 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c242
*+ bl_0_242 br_0_242 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c242
*+ bl_0_242 br_0_242 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c242
*+ bl_0_242 br_0_242 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c242
*+ bl_0_242 br_0_242 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c242
*+ bl_0_242 br_0_242 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c242
*+ bl_0_242 br_0_242 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c242
*+ bl_0_242 br_0_242 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c242
*+ bl_0_242 br_0_242 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c242
*+ bl_0_242 br_0_242 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c242
*+ bl_0_242 br_0_242 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c242
*+ bl_0_242 br_0_242 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c242
*+ bl_0_242 br_0_242 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c242
*+ bl_0_242 br_0_242 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c242
*+ bl_0_242 br_0_242 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c242
*+ bl_0_242 br_0_242 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c242
*+ bl_0_242 br_0_242 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c242
*+ bl_0_242 br_0_242 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c242
*+ bl_0_242 br_0_242 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c242
*+ bl_0_242 br_0_242 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c242
*+ bl_0_242 br_0_242 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c242
*+ bl_0_242 br_0_242 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c242
*+ bl_0_242 br_0_242 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c242
*+ bl_0_242 br_0_242 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c242
*+ bl_0_242 br_0_242 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c242
*+ bl_0_242 br_0_242 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c242
*+ bl_0_242 br_0_242 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c242
*+ bl_0_242 br_0_242 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c242
*+ bl_0_242 br_0_242 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c242
*+ bl_0_242 br_0_242 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c242
*+ bl_0_242 br_0_242 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c242
*+ bl_0_242 br_0_242 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c242
*+ bl_0_242 br_0_242 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c242
*+ bl_0_242 br_0_242 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c242
*+ bl_0_242 br_0_242 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c242
*+ bl_0_242 br_0_242 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c242
*+ bl_0_242 br_0_242 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c242
*+ bl_0_242 br_0_242 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c242
*+ bl_0_242 br_0_242 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c242
*+ bl_0_242 br_0_242 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c242
*+ bl_0_242 br_0_242 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c242
*+ bl_0_242 br_0_242 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c242
*+ bl_0_242 br_0_242 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c242
*+ bl_0_242 br_0_242 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c242
*+ bl_0_242 br_0_242 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c242
*+ bl_0_242 br_0_242 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c242
*+ bl_0_242 br_0_242 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c242
*+ bl_0_242 br_0_242 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c242
*+ bl_0_242 br_0_242 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c242
*+ bl_0_242 br_0_242 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c242
*+ bl_0_242 br_0_242 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c242
*+ bl_0_242 br_0_242 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c242
*+ bl_0_242 br_0_242 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c242
*+ bl_0_242 br_0_242 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c242
*+ bl_0_242 br_0_242 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c242
*+ bl_0_242 br_0_242 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c242
*+ bl_0_242 br_0_242 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c242
*+ bl_0_242 br_0_242 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c242
*+ bl_0_242 br_0_242 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c242
*+ bl_0_242 br_0_242 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c242
*+ bl_0_242 br_0_242 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c242
*+ bl_0_242 br_0_242 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c242
*+ bl_0_242 br_0_242 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c242
*+ bl_0_242 br_0_242 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c242
*+ bl_0_242 br_0_242 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c242
*+ bl_0_242 br_0_242 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c242
*+ bl_0_242 br_0_242 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c242
*+ bl_0_242 br_0_242 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c242
*+ bl_0_242 br_0_242 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c242
*+ bl_0_242 br_0_242 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c242
*+ bl_0_242 br_0_242 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c242
*+ bl_0_242 br_0_242 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c242
*+ bl_0_242 br_0_242 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c242
*+ bl_0_242 br_0_242 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c242
*+ bl_0_242 br_0_242 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c242
*+ bl_0_242 br_0_242 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c242
*+ bl_0_242 br_0_242 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c242
*+ bl_0_242 br_0_242 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c242
*+ bl_0_242 br_0_242 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c242
*+ bl_0_242 br_0_242 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c242
*+ bl_0_242 br_0_242 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c242
*+ bl_0_242 br_0_242 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c242
*+ bl_0_242 br_0_242 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c242
*+ bl_0_242 br_0_242 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c242
*+ bl_0_242 br_0_242 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c242
*+ bl_0_242 br_0_242 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c242
*+ bl_0_242 br_0_242 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c242
*+ bl_0_242 br_0_242 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c242
*+ bl_0_242 br_0_242 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c242
*+ bl_0_242 br_0_242 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c242
*+ bl_0_242 br_0_242 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c242
*+ bl_0_242 br_0_242 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c242
*+ bl_0_242 br_0_242 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c242
*+ bl_0_242 br_0_242 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c242
*+ bl_0_242 br_0_242 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c242
*+ bl_0_242 br_0_242 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c242
*+ bl_0_242 br_0_242 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c242
*+ bl_0_242 br_0_242 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c242
*+ bl_0_242 br_0_242 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c242
*+ bl_0_242 br_0_242 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c242
*+ bl_0_242 br_0_242 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c242
*+ bl_0_242 br_0_242 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c242
*+ bl_0_242 br_0_242 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c242
*+ bl_0_242 br_0_242 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c242
*+ bl_0_242 br_0_242 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c242
*+ bl_0_242 br_0_242 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c242
*+ bl_0_242 br_0_242 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c242
*+ bl_0_242 br_0_242 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c242
*+ bl_0_242 br_0_242 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c242
*+ bl_0_242 br_0_242 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c242
*+ bl_0_242 br_0_242 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c242
*+ bl_0_242 br_0_242 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c242
*+ bl_0_242 br_0_242 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c242
*+ bl_0_242 br_0_242 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c242
*+ bl_0_242 br_0_242 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c242
*+ bl_0_242 br_0_242 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c242
*+ bl_0_242 br_0_242 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c242
*+ bl_0_242 br_0_242 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c242
*+ bl_0_242 br_0_242 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c242
*+ bl_0_242 br_0_242 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c242
*+ bl_0_242 br_0_242 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c242
*+ bl_0_242 br_0_242 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c242
*+ bl_0_242 br_0_242 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c242
+ bl_0_242 br_0_242 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c243
+ bl_0_243 br_0_243 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c243
*+ bl_0_243 br_0_243 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c243
*+ bl_0_243 br_0_243 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c243
*+ bl_0_243 br_0_243 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c243
*+ bl_0_243 br_0_243 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c243
*+ bl_0_243 br_0_243 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c243
*+ bl_0_243 br_0_243 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c243
*+ bl_0_243 br_0_243 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c243
*+ bl_0_243 br_0_243 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c243
*+ bl_0_243 br_0_243 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c243
*+ bl_0_243 br_0_243 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c243
*+ bl_0_243 br_0_243 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c243
*+ bl_0_243 br_0_243 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c243
*+ bl_0_243 br_0_243 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c243
*+ bl_0_243 br_0_243 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c243
*+ bl_0_243 br_0_243 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c243
*+ bl_0_243 br_0_243 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c243
*+ bl_0_243 br_0_243 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c243
*+ bl_0_243 br_0_243 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c243
*+ bl_0_243 br_0_243 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c243
*+ bl_0_243 br_0_243 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c243
*+ bl_0_243 br_0_243 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c243
*+ bl_0_243 br_0_243 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c243
*+ bl_0_243 br_0_243 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c243
*+ bl_0_243 br_0_243 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c243
*+ bl_0_243 br_0_243 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c243
*+ bl_0_243 br_0_243 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c243
*+ bl_0_243 br_0_243 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c243
*+ bl_0_243 br_0_243 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c243
*+ bl_0_243 br_0_243 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c243
*+ bl_0_243 br_0_243 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c243
*+ bl_0_243 br_0_243 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c243
*+ bl_0_243 br_0_243 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c243
*+ bl_0_243 br_0_243 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c243
*+ bl_0_243 br_0_243 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c243
*+ bl_0_243 br_0_243 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c243
*+ bl_0_243 br_0_243 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c243
*+ bl_0_243 br_0_243 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c243
*+ bl_0_243 br_0_243 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c243
*+ bl_0_243 br_0_243 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c243
*+ bl_0_243 br_0_243 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c243
*+ bl_0_243 br_0_243 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c243
*+ bl_0_243 br_0_243 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c243
*+ bl_0_243 br_0_243 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c243
*+ bl_0_243 br_0_243 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c243
*+ bl_0_243 br_0_243 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c243
*+ bl_0_243 br_0_243 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c243
*+ bl_0_243 br_0_243 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c243
*+ bl_0_243 br_0_243 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c243
*+ bl_0_243 br_0_243 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c243
*+ bl_0_243 br_0_243 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c243
*+ bl_0_243 br_0_243 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c243
*+ bl_0_243 br_0_243 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c243
*+ bl_0_243 br_0_243 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c243
*+ bl_0_243 br_0_243 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c243
*+ bl_0_243 br_0_243 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c243
*+ bl_0_243 br_0_243 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c243
*+ bl_0_243 br_0_243 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c243
*+ bl_0_243 br_0_243 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c243
*+ bl_0_243 br_0_243 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c243
*+ bl_0_243 br_0_243 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c243
*+ bl_0_243 br_0_243 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c243
*+ bl_0_243 br_0_243 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c243
*+ bl_0_243 br_0_243 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c243
*+ bl_0_243 br_0_243 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c243
*+ bl_0_243 br_0_243 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c243
*+ bl_0_243 br_0_243 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c243
*+ bl_0_243 br_0_243 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c243
*+ bl_0_243 br_0_243 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c243
*+ bl_0_243 br_0_243 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c243
*+ bl_0_243 br_0_243 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c243
*+ bl_0_243 br_0_243 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c243
*+ bl_0_243 br_0_243 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c243
*+ bl_0_243 br_0_243 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c243
*+ bl_0_243 br_0_243 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c243
*+ bl_0_243 br_0_243 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c243
*+ bl_0_243 br_0_243 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c243
*+ bl_0_243 br_0_243 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c243
*+ bl_0_243 br_0_243 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c243
*+ bl_0_243 br_0_243 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c243
*+ bl_0_243 br_0_243 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c243
*+ bl_0_243 br_0_243 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c243
*+ bl_0_243 br_0_243 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c243
*+ bl_0_243 br_0_243 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c243
*+ bl_0_243 br_0_243 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c243
*+ bl_0_243 br_0_243 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c243
*+ bl_0_243 br_0_243 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c243
*+ bl_0_243 br_0_243 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c243
*+ bl_0_243 br_0_243 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c243
*+ bl_0_243 br_0_243 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c243
*+ bl_0_243 br_0_243 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c243
*+ bl_0_243 br_0_243 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c243
*+ bl_0_243 br_0_243 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c243
*+ bl_0_243 br_0_243 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c243
*+ bl_0_243 br_0_243 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c243
*+ bl_0_243 br_0_243 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c243
*+ bl_0_243 br_0_243 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c243
*+ bl_0_243 br_0_243 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c243
*+ bl_0_243 br_0_243 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c243
*+ bl_0_243 br_0_243 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c243
*+ bl_0_243 br_0_243 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c243
*+ bl_0_243 br_0_243 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c243
*+ bl_0_243 br_0_243 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c243
*+ bl_0_243 br_0_243 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c243
*+ bl_0_243 br_0_243 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c243
*+ bl_0_243 br_0_243 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c243
*+ bl_0_243 br_0_243 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c243
*+ bl_0_243 br_0_243 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c243
*+ bl_0_243 br_0_243 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c243
*+ bl_0_243 br_0_243 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c243
*+ bl_0_243 br_0_243 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c243
*+ bl_0_243 br_0_243 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c243
*+ bl_0_243 br_0_243 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c243
*+ bl_0_243 br_0_243 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c243
*+ bl_0_243 br_0_243 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c243
*+ bl_0_243 br_0_243 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c243
*+ bl_0_243 br_0_243 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c243
*+ bl_0_243 br_0_243 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c243
*+ bl_0_243 br_0_243 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c243
*+ bl_0_243 br_0_243 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c243
*+ bl_0_243 br_0_243 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c243
*+ bl_0_243 br_0_243 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c243
*+ bl_0_243 br_0_243 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c243
*+ bl_0_243 br_0_243 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c243
*+ bl_0_243 br_0_243 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c243
*+ bl_0_243 br_0_243 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c243
*+ bl_0_243 br_0_243 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c243
+ bl_0_243 br_0_243 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c244
+ bl_0_244 br_0_244 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c244
*+ bl_0_244 br_0_244 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c244
*+ bl_0_244 br_0_244 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c244
*+ bl_0_244 br_0_244 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c244
*+ bl_0_244 br_0_244 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c244
*+ bl_0_244 br_0_244 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c244
*+ bl_0_244 br_0_244 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c244
*+ bl_0_244 br_0_244 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c244
*+ bl_0_244 br_0_244 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c244
*+ bl_0_244 br_0_244 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c244
*+ bl_0_244 br_0_244 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c244
*+ bl_0_244 br_0_244 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c244
*+ bl_0_244 br_0_244 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c244
*+ bl_0_244 br_0_244 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c244
*+ bl_0_244 br_0_244 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c244
*+ bl_0_244 br_0_244 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c244
*+ bl_0_244 br_0_244 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c244
*+ bl_0_244 br_0_244 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c244
*+ bl_0_244 br_0_244 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c244
*+ bl_0_244 br_0_244 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c244
*+ bl_0_244 br_0_244 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c244
*+ bl_0_244 br_0_244 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c244
*+ bl_0_244 br_0_244 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c244
*+ bl_0_244 br_0_244 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c244
*+ bl_0_244 br_0_244 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c244
*+ bl_0_244 br_0_244 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c244
*+ bl_0_244 br_0_244 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c244
*+ bl_0_244 br_0_244 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c244
*+ bl_0_244 br_0_244 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c244
*+ bl_0_244 br_0_244 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c244
*+ bl_0_244 br_0_244 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c244
*+ bl_0_244 br_0_244 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c244
*+ bl_0_244 br_0_244 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c244
*+ bl_0_244 br_0_244 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c244
*+ bl_0_244 br_0_244 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c244
*+ bl_0_244 br_0_244 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c244
*+ bl_0_244 br_0_244 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c244
*+ bl_0_244 br_0_244 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c244
*+ bl_0_244 br_0_244 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c244
*+ bl_0_244 br_0_244 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c244
*+ bl_0_244 br_0_244 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c244
*+ bl_0_244 br_0_244 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c244
*+ bl_0_244 br_0_244 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c244
*+ bl_0_244 br_0_244 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c244
*+ bl_0_244 br_0_244 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c244
*+ bl_0_244 br_0_244 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c244
*+ bl_0_244 br_0_244 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c244
*+ bl_0_244 br_0_244 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c244
*+ bl_0_244 br_0_244 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c244
*+ bl_0_244 br_0_244 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c244
*+ bl_0_244 br_0_244 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c244
*+ bl_0_244 br_0_244 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c244
*+ bl_0_244 br_0_244 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c244
*+ bl_0_244 br_0_244 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c244
*+ bl_0_244 br_0_244 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c244
*+ bl_0_244 br_0_244 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c244
*+ bl_0_244 br_0_244 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c244
*+ bl_0_244 br_0_244 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c244
*+ bl_0_244 br_0_244 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c244
*+ bl_0_244 br_0_244 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c244
*+ bl_0_244 br_0_244 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c244
*+ bl_0_244 br_0_244 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c244
*+ bl_0_244 br_0_244 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c244
*+ bl_0_244 br_0_244 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c244
*+ bl_0_244 br_0_244 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c244
*+ bl_0_244 br_0_244 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c244
*+ bl_0_244 br_0_244 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c244
*+ bl_0_244 br_0_244 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c244
*+ bl_0_244 br_0_244 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c244
*+ bl_0_244 br_0_244 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c244
*+ bl_0_244 br_0_244 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c244
*+ bl_0_244 br_0_244 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c244
*+ bl_0_244 br_0_244 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c244
*+ bl_0_244 br_0_244 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c244
*+ bl_0_244 br_0_244 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c244
*+ bl_0_244 br_0_244 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c244
*+ bl_0_244 br_0_244 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c244
*+ bl_0_244 br_0_244 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c244
*+ bl_0_244 br_0_244 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c244
*+ bl_0_244 br_0_244 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c244
*+ bl_0_244 br_0_244 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c244
*+ bl_0_244 br_0_244 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c244
*+ bl_0_244 br_0_244 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c244
*+ bl_0_244 br_0_244 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c244
*+ bl_0_244 br_0_244 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c244
*+ bl_0_244 br_0_244 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c244
*+ bl_0_244 br_0_244 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c244
*+ bl_0_244 br_0_244 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c244
*+ bl_0_244 br_0_244 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c244
*+ bl_0_244 br_0_244 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c244
*+ bl_0_244 br_0_244 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c244
*+ bl_0_244 br_0_244 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c244
*+ bl_0_244 br_0_244 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c244
*+ bl_0_244 br_0_244 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c244
*+ bl_0_244 br_0_244 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c244
*+ bl_0_244 br_0_244 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c244
*+ bl_0_244 br_0_244 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c244
*+ bl_0_244 br_0_244 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c244
*+ bl_0_244 br_0_244 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c244
*+ bl_0_244 br_0_244 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c244
*+ bl_0_244 br_0_244 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c244
*+ bl_0_244 br_0_244 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c244
*+ bl_0_244 br_0_244 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c244
*+ bl_0_244 br_0_244 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c244
*+ bl_0_244 br_0_244 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c244
*+ bl_0_244 br_0_244 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c244
*+ bl_0_244 br_0_244 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c244
*+ bl_0_244 br_0_244 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c244
*+ bl_0_244 br_0_244 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c244
*+ bl_0_244 br_0_244 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c244
*+ bl_0_244 br_0_244 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c244
*+ bl_0_244 br_0_244 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c244
*+ bl_0_244 br_0_244 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c244
*+ bl_0_244 br_0_244 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c244
*+ bl_0_244 br_0_244 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c244
*+ bl_0_244 br_0_244 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c244
*+ bl_0_244 br_0_244 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c244
*+ bl_0_244 br_0_244 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c244
*+ bl_0_244 br_0_244 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c244
*+ bl_0_244 br_0_244 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c244
*+ bl_0_244 br_0_244 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c244
*+ bl_0_244 br_0_244 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c244
*+ bl_0_244 br_0_244 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c244
*+ bl_0_244 br_0_244 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c244
*+ bl_0_244 br_0_244 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c244
*+ bl_0_244 br_0_244 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c244
*+ bl_0_244 br_0_244 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c244
+ bl_0_244 br_0_244 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c245
+ bl_0_245 br_0_245 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c245
*+ bl_0_245 br_0_245 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c245
*+ bl_0_245 br_0_245 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c245
*+ bl_0_245 br_0_245 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c245
*+ bl_0_245 br_0_245 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c245
*+ bl_0_245 br_0_245 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c245
*+ bl_0_245 br_0_245 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c245
*+ bl_0_245 br_0_245 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c245
*+ bl_0_245 br_0_245 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c245
*+ bl_0_245 br_0_245 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c245
*+ bl_0_245 br_0_245 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c245
*+ bl_0_245 br_0_245 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c245
*+ bl_0_245 br_0_245 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c245
*+ bl_0_245 br_0_245 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c245
*+ bl_0_245 br_0_245 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c245
*+ bl_0_245 br_0_245 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c245
*+ bl_0_245 br_0_245 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c245
*+ bl_0_245 br_0_245 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c245
*+ bl_0_245 br_0_245 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c245
*+ bl_0_245 br_0_245 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c245
*+ bl_0_245 br_0_245 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c245
*+ bl_0_245 br_0_245 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c245
*+ bl_0_245 br_0_245 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c245
*+ bl_0_245 br_0_245 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c245
*+ bl_0_245 br_0_245 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c245
*+ bl_0_245 br_0_245 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c245
*+ bl_0_245 br_0_245 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c245
*+ bl_0_245 br_0_245 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c245
*+ bl_0_245 br_0_245 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c245
*+ bl_0_245 br_0_245 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c245
*+ bl_0_245 br_0_245 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c245
*+ bl_0_245 br_0_245 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c245
*+ bl_0_245 br_0_245 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c245
*+ bl_0_245 br_0_245 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c245
*+ bl_0_245 br_0_245 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c245
*+ bl_0_245 br_0_245 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c245
*+ bl_0_245 br_0_245 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c245
*+ bl_0_245 br_0_245 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c245
*+ bl_0_245 br_0_245 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c245
*+ bl_0_245 br_0_245 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c245
*+ bl_0_245 br_0_245 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c245
*+ bl_0_245 br_0_245 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c245
*+ bl_0_245 br_0_245 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c245
*+ bl_0_245 br_0_245 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c245
*+ bl_0_245 br_0_245 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c245
*+ bl_0_245 br_0_245 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c245
*+ bl_0_245 br_0_245 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c245
*+ bl_0_245 br_0_245 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c245
*+ bl_0_245 br_0_245 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c245
*+ bl_0_245 br_0_245 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c245
*+ bl_0_245 br_0_245 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c245
*+ bl_0_245 br_0_245 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c245
*+ bl_0_245 br_0_245 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c245
*+ bl_0_245 br_0_245 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c245
*+ bl_0_245 br_0_245 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c245
*+ bl_0_245 br_0_245 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c245
*+ bl_0_245 br_0_245 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c245
*+ bl_0_245 br_0_245 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c245
*+ bl_0_245 br_0_245 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c245
*+ bl_0_245 br_0_245 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c245
*+ bl_0_245 br_0_245 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c245
*+ bl_0_245 br_0_245 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c245
*+ bl_0_245 br_0_245 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c245
*+ bl_0_245 br_0_245 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c245
*+ bl_0_245 br_0_245 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c245
*+ bl_0_245 br_0_245 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c245
*+ bl_0_245 br_0_245 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c245
*+ bl_0_245 br_0_245 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c245
*+ bl_0_245 br_0_245 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c245
*+ bl_0_245 br_0_245 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c245
*+ bl_0_245 br_0_245 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c245
*+ bl_0_245 br_0_245 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c245
*+ bl_0_245 br_0_245 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c245
*+ bl_0_245 br_0_245 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c245
*+ bl_0_245 br_0_245 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c245
*+ bl_0_245 br_0_245 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c245
*+ bl_0_245 br_0_245 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c245
*+ bl_0_245 br_0_245 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c245
*+ bl_0_245 br_0_245 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c245
*+ bl_0_245 br_0_245 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c245
*+ bl_0_245 br_0_245 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c245
*+ bl_0_245 br_0_245 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c245
*+ bl_0_245 br_0_245 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c245
*+ bl_0_245 br_0_245 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c245
*+ bl_0_245 br_0_245 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c245
*+ bl_0_245 br_0_245 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c245
*+ bl_0_245 br_0_245 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c245
*+ bl_0_245 br_0_245 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c245
*+ bl_0_245 br_0_245 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c245
*+ bl_0_245 br_0_245 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c245
*+ bl_0_245 br_0_245 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c245
*+ bl_0_245 br_0_245 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c245
*+ bl_0_245 br_0_245 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c245
*+ bl_0_245 br_0_245 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c245
*+ bl_0_245 br_0_245 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c245
*+ bl_0_245 br_0_245 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c245
*+ bl_0_245 br_0_245 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c245
*+ bl_0_245 br_0_245 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c245
*+ bl_0_245 br_0_245 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c245
*+ bl_0_245 br_0_245 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c245
*+ bl_0_245 br_0_245 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c245
*+ bl_0_245 br_0_245 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c245
*+ bl_0_245 br_0_245 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c245
*+ bl_0_245 br_0_245 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c245
*+ bl_0_245 br_0_245 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c245
*+ bl_0_245 br_0_245 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c245
*+ bl_0_245 br_0_245 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c245
*+ bl_0_245 br_0_245 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c245
*+ bl_0_245 br_0_245 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c245
*+ bl_0_245 br_0_245 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c245
*+ bl_0_245 br_0_245 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c245
*+ bl_0_245 br_0_245 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c245
*+ bl_0_245 br_0_245 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c245
*+ bl_0_245 br_0_245 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c245
*+ bl_0_245 br_0_245 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c245
*+ bl_0_245 br_0_245 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c245
*+ bl_0_245 br_0_245 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c245
*+ bl_0_245 br_0_245 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c245
*+ bl_0_245 br_0_245 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c245
*+ bl_0_245 br_0_245 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c245
*+ bl_0_245 br_0_245 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c245
*+ bl_0_245 br_0_245 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c245
*+ bl_0_245 br_0_245 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c245
*+ bl_0_245 br_0_245 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c245
*+ bl_0_245 br_0_245 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c245
*+ bl_0_245 br_0_245 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c245
*+ bl_0_245 br_0_245 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c245
+ bl_0_245 br_0_245 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c246
+ bl_0_246 br_0_246 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c246
*+ bl_0_246 br_0_246 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c246
*+ bl_0_246 br_0_246 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c246
*+ bl_0_246 br_0_246 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c246
*+ bl_0_246 br_0_246 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c246
*+ bl_0_246 br_0_246 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c246
*+ bl_0_246 br_0_246 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c246
*+ bl_0_246 br_0_246 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c246
*+ bl_0_246 br_0_246 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c246
*+ bl_0_246 br_0_246 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c246
*+ bl_0_246 br_0_246 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c246
*+ bl_0_246 br_0_246 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c246
*+ bl_0_246 br_0_246 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c246
*+ bl_0_246 br_0_246 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c246
*+ bl_0_246 br_0_246 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c246
*+ bl_0_246 br_0_246 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c246
*+ bl_0_246 br_0_246 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c246
*+ bl_0_246 br_0_246 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c246
*+ bl_0_246 br_0_246 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c246
*+ bl_0_246 br_0_246 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c246
*+ bl_0_246 br_0_246 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c246
*+ bl_0_246 br_0_246 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c246
*+ bl_0_246 br_0_246 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c246
*+ bl_0_246 br_0_246 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c246
*+ bl_0_246 br_0_246 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c246
*+ bl_0_246 br_0_246 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c246
*+ bl_0_246 br_0_246 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c246
*+ bl_0_246 br_0_246 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c246
*+ bl_0_246 br_0_246 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c246
*+ bl_0_246 br_0_246 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c246
*+ bl_0_246 br_0_246 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c246
*+ bl_0_246 br_0_246 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c246
*+ bl_0_246 br_0_246 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c246
*+ bl_0_246 br_0_246 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c246
*+ bl_0_246 br_0_246 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c246
*+ bl_0_246 br_0_246 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c246
*+ bl_0_246 br_0_246 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c246
*+ bl_0_246 br_0_246 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c246
*+ bl_0_246 br_0_246 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c246
*+ bl_0_246 br_0_246 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c246
*+ bl_0_246 br_0_246 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c246
*+ bl_0_246 br_0_246 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c246
*+ bl_0_246 br_0_246 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c246
*+ bl_0_246 br_0_246 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c246
*+ bl_0_246 br_0_246 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c246
*+ bl_0_246 br_0_246 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c246
*+ bl_0_246 br_0_246 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c246
*+ bl_0_246 br_0_246 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c246
*+ bl_0_246 br_0_246 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c246
*+ bl_0_246 br_0_246 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c246
*+ bl_0_246 br_0_246 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c246
*+ bl_0_246 br_0_246 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c246
*+ bl_0_246 br_0_246 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c246
*+ bl_0_246 br_0_246 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c246
*+ bl_0_246 br_0_246 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c246
*+ bl_0_246 br_0_246 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c246
*+ bl_0_246 br_0_246 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c246
*+ bl_0_246 br_0_246 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c246
*+ bl_0_246 br_0_246 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c246
*+ bl_0_246 br_0_246 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c246
*+ bl_0_246 br_0_246 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c246
*+ bl_0_246 br_0_246 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c246
*+ bl_0_246 br_0_246 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c246
*+ bl_0_246 br_0_246 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c246
*+ bl_0_246 br_0_246 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c246
*+ bl_0_246 br_0_246 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c246
*+ bl_0_246 br_0_246 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c246
*+ bl_0_246 br_0_246 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c246
*+ bl_0_246 br_0_246 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c246
*+ bl_0_246 br_0_246 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c246
*+ bl_0_246 br_0_246 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c246
*+ bl_0_246 br_0_246 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c246
*+ bl_0_246 br_0_246 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c246
*+ bl_0_246 br_0_246 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c246
*+ bl_0_246 br_0_246 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c246
*+ bl_0_246 br_0_246 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c246
*+ bl_0_246 br_0_246 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c246
*+ bl_0_246 br_0_246 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c246
*+ bl_0_246 br_0_246 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c246
*+ bl_0_246 br_0_246 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c246
*+ bl_0_246 br_0_246 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c246
*+ bl_0_246 br_0_246 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c246
*+ bl_0_246 br_0_246 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c246
*+ bl_0_246 br_0_246 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c246
*+ bl_0_246 br_0_246 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c246
*+ bl_0_246 br_0_246 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c246
*+ bl_0_246 br_0_246 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c246
*+ bl_0_246 br_0_246 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c246
*+ bl_0_246 br_0_246 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c246
*+ bl_0_246 br_0_246 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c246
*+ bl_0_246 br_0_246 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c246
*+ bl_0_246 br_0_246 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c246
*+ bl_0_246 br_0_246 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c246
*+ bl_0_246 br_0_246 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c246
*+ bl_0_246 br_0_246 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c246
*+ bl_0_246 br_0_246 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c246
*+ bl_0_246 br_0_246 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c246
*+ bl_0_246 br_0_246 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c246
*+ bl_0_246 br_0_246 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c246
*+ bl_0_246 br_0_246 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c246
*+ bl_0_246 br_0_246 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c246
*+ bl_0_246 br_0_246 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c246
*+ bl_0_246 br_0_246 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c246
*+ bl_0_246 br_0_246 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c246
*+ bl_0_246 br_0_246 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c246
*+ bl_0_246 br_0_246 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c246
*+ bl_0_246 br_0_246 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c246
*+ bl_0_246 br_0_246 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c246
*+ bl_0_246 br_0_246 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c246
*+ bl_0_246 br_0_246 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c246
*+ bl_0_246 br_0_246 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c246
*+ bl_0_246 br_0_246 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c246
*+ bl_0_246 br_0_246 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c246
*+ bl_0_246 br_0_246 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c246
*+ bl_0_246 br_0_246 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c246
*+ bl_0_246 br_0_246 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c246
*+ bl_0_246 br_0_246 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c246
*+ bl_0_246 br_0_246 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c246
*+ bl_0_246 br_0_246 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c246
*+ bl_0_246 br_0_246 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c246
*+ bl_0_246 br_0_246 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c246
*+ bl_0_246 br_0_246 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c246
*+ bl_0_246 br_0_246 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c246
*+ bl_0_246 br_0_246 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c246
*+ bl_0_246 br_0_246 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c246
*+ bl_0_246 br_0_246 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c246
*+ bl_0_246 br_0_246 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c246
+ bl_0_246 br_0_246 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c247
+ bl_0_247 br_0_247 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c247
*+ bl_0_247 br_0_247 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c247
*+ bl_0_247 br_0_247 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c247
*+ bl_0_247 br_0_247 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c247
*+ bl_0_247 br_0_247 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c247
*+ bl_0_247 br_0_247 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c247
*+ bl_0_247 br_0_247 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c247
*+ bl_0_247 br_0_247 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c247
*+ bl_0_247 br_0_247 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c247
*+ bl_0_247 br_0_247 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c247
*+ bl_0_247 br_0_247 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c247
*+ bl_0_247 br_0_247 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c247
*+ bl_0_247 br_0_247 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c247
*+ bl_0_247 br_0_247 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c247
*+ bl_0_247 br_0_247 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c247
*+ bl_0_247 br_0_247 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c247
*+ bl_0_247 br_0_247 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c247
*+ bl_0_247 br_0_247 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c247
*+ bl_0_247 br_0_247 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c247
*+ bl_0_247 br_0_247 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c247
*+ bl_0_247 br_0_247 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c247
*+ bl_0_247 br_0_247 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c247
*+ bl_0_247 br_0_247 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c247
*+ bl_0_247 br_0_247 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c247
*+ bl_0_247 br_0_247 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c247
*+ bl_0_247 br_0_247 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c247
*+ bl_0_247 br_0_247 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c247
*+ bl_0_247 br_0_247 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c247
*+ bl_0_247 br_0_247 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c247
*+ bl_0_247 br_0_247 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c247
*+ bl_0_247 br_0_247 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c247
*+ bl_0_247 br_0_247 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c247
*+ bl_0_247 br_0_247 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c247
*+ bl_0_247 br_0_247 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c247
*+ bl_0_247 br_0_247 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c247
*+ bl_0_247 br_0_247 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c247
*+ bl_0_247 br_0_247 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c247
*+ bl_0_247 br_0_247 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c247
*+ bl_0_247 br_0_247 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c247
*+ bl_0_247 br_0_247 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c247
*+ bl_0_247 br_0_247 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c247
*+ bl_0_247 br_0_247 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c247
*+ bl_0_247 br_0_247 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c247
*+ bl_0_247 br_0_247 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c247
*+ bl_0_247 br_0_247 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c247
*+ bl_0_247 br_0_247 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c247
*+ bl_0_247 br_0_247 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c247
*+ bl_0_247 br_0_247 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c247
*+ bl_0_247 br_0_247 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c247
*+ bl_0_247 br_0_247 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c247
*+ bl_0_247 br_0_247 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c247
*+ bl_0_247 br_0_247 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c247
*+ bl_0_247 br_0_247 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c247
*+ bl_0_247 br_0_247 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c247
*+ bl_0_247 br_0_247 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c247
*+ bl_0_247 br_0_247 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c247
*+ bl_0_247 br_0_247 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c247
*+ bl_0_247 br_0_247 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c247
*+ bl_0_247 br_0_247 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c247
*+ bl_0_247 br_0_247 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c247
*+ bl_0_247 br_0_247 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c247
*+ bl_0_247 br_0_247 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c247
*+ bl_0_247 br_0_247 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c247
*+ bl_0_247 br_0_247 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c247
*+ bl_0_247 br_0_247 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c247
*+ bl_0_247 br_0_247 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c247
*+ bl_0_247 br_0_247 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c247
*+ bl_0_247 br_0_247 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c247
*+ bl_0_247 br_0_247 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c247
*+ bl_0_247 br_0_247 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c247
*+ bl_0_247 br_0_247 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c247
*+ bl_0_247 br_0_247 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c247
*+ bl_0_247 br_0_247 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c247
*+ bl_0_247 br_0_247 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c247
*+ bl_0_247 br_0_247 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c247
*+ bl_0_247 br_0_247 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c247
*+ bl_0_247 br_0_247 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c247
*+ bl_0_247 br_0_247 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c247
*+ bl_0_247 br_0_247 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c247
*+ bl_0_247 br_0_247 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c247
*+ bl_0_247 br_0_247 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c247
*+ bl_0_247 br_0_247 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c247
*+ bl_0_247 br_0_247 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c247
*+ bl_0_247 br_0_247 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c247
*+ bl_0_247 br_0_247 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c247
*+ bl_0_247 br_0_247 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c247
*+ bl_0_247 br_0_247 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c247
*+ bl_0_247 br_0_247 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c247
*+ bl_0_247 br_0_247 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c247
*+ bl_0_247 br_0_247 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c247
*+ bl_0_247 br_0_247 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c247
*+ bl_0_247 br_0_247 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c247
*+ bl_0_247 br_0_247 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c247
*+ bl_0_247 br_0_247 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c247
*+ bl_0_247 br_0_247 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c247
*+ bl_0_247 br_0_247 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c247
*+ bl_0_247 br_0_247 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c247
*+ bl_0_247 br_0_247 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c247
*+ bl_0_247 br_0_247 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c247
*+ bl_0_247 br_0_247 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c247
*+ bl_0_247 br_0_247 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c247
*+ bl_0_247 br_0_247 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c247
*+ bl_0_247 br_0_247 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c247
*+ bl_0_247 br_0_247 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c247
*+ bl_0_247 br_0_247 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c247
*+ bl_0_247 br_0_247 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c247
*+ bl_0_247 br_0_247 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c247
*+ bl_0_247 br_0_247 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c247
*+ bl_0_247 br_0_247 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c247
*+ bl_0_247 br_0_247 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c247
*+ bl_0_247 br_0_247 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c247
*+ bl_0_247 br_0_247 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c247
*+ bl_0_247 br_0_247 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c247
*+ bl_0_247 br_0_247 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c247
*+ bl_0_247 br_0_247 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c247
*+ bl_0_247 br_0_247 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c247
*+ bl_0_247 br_0_247 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c247
*+ bl_0_247 br_0_247 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c247
*+ bl_0_247 br_0_247 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c247
*+ bl_0_247 br_0_247 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c247
*+ bl_0_247 br_0_247 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c247
*+ bl_0_247 br_0_247 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c247
*+ bl_0_247 br_0_247 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c247
*+ bl_0_247 br_0_247 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c247
*+ bl_0_247 br_0_247 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c247
*+ bl_0_247 br_0_247 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c247
*+ bl_0_247 br_0_247 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c247
+ bl_0_247 br_0_247 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c248
+ bl_0_248 br_0_248 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c248
*+ bl_0_248 br_0_248 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c248
*+ bl_0_248 br_0_248 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c248
*+ bl_0_248 br_0_248 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c248
*+ bl_0_248 br_0_248 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c248
*+ bl_0_248 br_0_248 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c248
*+ bl_0_248 br_0_248 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c248
*+ bl_0_248 br_0_248 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c248
*+ bl_0_248 br_0_248 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c248
*+ bl_0_248 br_0_248 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c248
*+ bl_0_248 br_0_248 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c248
*+ bl_0_248 br_0_248 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c248
*+ bl_0_248 br_0_248 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c248
*+ bl_0_248 br_0_248 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c248
*+ bl_0_248 br_0_248 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c248
*+ bl_0_248 br_0_248 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c248
*+ bl_0_248 br_0_248 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c248
*+ bl_0_248 br_0_248 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c248
*+ bl_0_248 br_0_248 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c248
*+ bl_0_248 br_0_248 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c248
*+ bl_0_248 br_0_248 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c248
*+ bl_0_248 br_0_248 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c248
*+ bl_0_248 br_0_248 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c248
*+ bl_0_248 br_0_248 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c248
*+ bl_0_248 br_0_248 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c248
*+ bl_0_248 br_0_248 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c248
*+ bl_0_248 br_0_248 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c248
*+ bl_0_248 br_0_248 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c248
*+ bl_0_248 br_0_248 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c248
*+ bl_0_248 br_0_248 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c248
*+ bl_0_248 br_0_248 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c248
*+ bl_0_248 br_0_248 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c248
*+ bl_0_248 br_0_248 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c248
*+ bl_0_248 br_0_248 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c248
*+ bl_0_248 br_0_248 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c248
*+ bl_0_248 br_0_248 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c248
*+ bl_0_248 br_0_248 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c248
*+ bl_0_248 br_0_248 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c248
*+ bl_0_248 br_0_248 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c248
*+ bl_0_248 br_0_248 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c248
*+ bl_0_248 br_0_248 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c248
*+ bl_0_248 br_0_248 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c248
*+ bl_0_248 br_0_248 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c248
*+ bl_0_248 br_0_248 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c248
*+ bl_0_248 br_0_248 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c248
*+ bl_0_248 br_0_248 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c248
*+ bl_0_248 br_0_248 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c248
*+ bl_0_248 br_0_248 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c248
*+ bl_0_248 br_0_248 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c248
*+ bl_0_248 br_0_248 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c248
*+ bl_0_248 br_0_248 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c248
*+ bl_0_248 br_0_248 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c248
*+ bl_0_248 br_0_248 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c248
*+ bl_0_248 br_0_248 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c248
*+ bl_0_248 br_0_248 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c248
*+ bl_0_248 br_0_248 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c248
*+ bl_0_248 br_0_248 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c248
*+ bl_0_248 br_0_248 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c248
*+ bl_0_248 br_0_248 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c248
*+ bl_0_248 br_0_248 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c248
*+ bl_0_248 br_0_248 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c248
*+ bl_0_248 br_0_248 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c248
*+ bl_0_248 br_0_248 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c248
*+ bl_0_248 br_0_248 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c248
*+ bl_0_248 br_0_248 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c248
*+ bl_0_248 br_0_248 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c248
*+ bl_0_248 br_0_248 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c248
*+ bl_0_248 br_0_248 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c248
*+ bl_0_248 br_0_248 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c248
*+ bl_0_248 br_0_248 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c248
*+ bl_0_248 br_0_248 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c248
*+ bl_0_248 br_0_248 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c248
*+ bl_0_248 br_0_248 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c248
*+ bl_0_248 br_0_248 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c248
*+ bl_0_248 br_0_248 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c248
*+ bl_0_248 br_0_248 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c248
*+ bl_0_248 br_0_248 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c248
*+ bl_0_248 br_0_248 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c248
*+ bl_0_248 br_0_248 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c248
*+ bl_0_248 br_0_248 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c248
*+ bl_0_248 br_0_248 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c248
*+ bl_0_248 br_0_248 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c248
*+ bl_0_248 br_0_248 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c248
*+ bl_0_248 br_0_248 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c248
*+ bl_0_248 br_0_248 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c248
*+ bl_0_248 br_0_248 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c248
*+ bl_0_248 br_0_248 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c248
*+ bl_0_248 br_0_248 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c248
*+ bl_0_248 br_0_248 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c248
*+ bl_0_248 br_0_248 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c248
*+ bl_0_248 br_0_248 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c248
*+ bl_0_248 br_0_248 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c248
*+ bl_0_248 br_0_248 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c248
*+ bl_0_248 br_0_248 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c248
*+ bl_0_248 br_0_248 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c248
*+ bl_0_248 br_0_248 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c248
*+ bl_0_248 br_0_248 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c248
*+ bl_0_248 br_0_248 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c248
*+ bl_0_248 br_0_248 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c248
*+ bl_0_248 br_0_248 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c248
*+ bl_0_248 br_0_248 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c248
*+ bl_0_248 br_0_248 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c248
*+ bl_0_248 br_0_248 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c248
*+ bl_0_248 br_0_248 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c248
*+ bl_0_248 br_0_248 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c248
*+ bl_0_248 br_0_248 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c248
*+ bl_0_248 br_0_248 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c248
*+ bl_0_248 br_0_248 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c248
*+ bl_0_248 br_0_248 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c248
*+ bl_0_248 br_0_248 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c248
*+ bl_0_248 br_0_248 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c248
*+ bl_0_248 br_0_248 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c248
*+ bl_0_248 br_0_248 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c248
*+ bl_0_248 br_0_248 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c248
*+ bl_0_248 br_0_248 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c248
*+ bl_0_248 br_0_248 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c248
*+ bl_0_248 br_0_248 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c248
*+ bl_0_248 br_0_248 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c248
*+ bl_0_248 br_0_248 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c248
*+ bl_0_248 br_0_248 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c248
*+ bl_0_248 br_0_248 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c248
*+ bl_0_248 br_0_248 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c248
*+ bl_0_248 br_0_248 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c248
*+ bl_0_248 br_0_248 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c248
*+ bl_0_248 br_0_248 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c248
*+ bl_0_248 br_0_248 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c248
*+ bl_0_248 br_0_248 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c248
+ bl_0_248 br_0_248 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c249
+ bl_0_249 br_0_249 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c249
*+ bl_0_249 br_0_249 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c249
*+ bl_0_249 br_0_249 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c249
*+ bl_0_249 br_0_249 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c249
*+ bl_0_249 br_0_249 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c249
*+ bl_0_249 br_0_249 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c249
*+ bl_0_249 br_0_249 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c249
*+ bl_0_249 br_0_249 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c249
*+ bl_0_249 br_0_249 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c249
*+ bl_0_249 br_0_249 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c249
*+ bl_0_249 br_0_249 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c249
*+ bl_0_249 br_0_249 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c249
*+ bl_0_249 br_0_249 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c249
*+ bl_0_249 br_0_249 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c249
*+ bl_0_249 br_0_249 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c249
*+ bl_0_249 br_0_249 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c249
*+ bl_0_249 br_0_249 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c249
*+ bl_0_249 br_0_249 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c249
*+ bl_0_249 br_0_249 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c249
*+ bl_0_249 br_0_249 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c249
*+ bl_0_249 br_0_249 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c249
*+ bl_0_249 br_0_249 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c249
*+ bl_0_249 br_0_249 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c249
*+ bl_0_249 br_0_249 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c249
*+ bl_0_249 br_0_249 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c249
*+ bl_0_249 br_0_249 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c249
*+ bl_0_249 br_0_249 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c249
*+ bl_0_249 br_0_249 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c249
*+ bl_0_249 br_0_249 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c249
*+ bl_0_249 br_0_249 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c249
*+ bl_0_249 br_0_249 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c249
*+ bl_0_249 br_0_249 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c249
*+ bl_0_249 br_0_249 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c249
*+ bl_0_249 br_0_249 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c249
*+ bl_0_249 br_0_249 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c249
*+ bl_0_249 br_0_249 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c249
*+ bl_0_249 br_0_249 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c249
*+ bl_0_249 br_0_249 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c249
*+ bl_0_249 br_0_249 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c249
*+ bl_0_249 br_0_249 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c249
*+ bl_0_249 br_0_249 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c249
*+ bl_0_249 br_0_249 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c249
*+ bl_0_249 br_0_249 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c249
*+ bl_0_249 br_0_249 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c249
*+ bl_0_249 br_0_249 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c249
*+ bl_0_249 br_0_249 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c249
*+ bl_0_249 br_0_249 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c249
*+ bl_0_249 br_0_249 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c249
*+ bl_0_249 br_0_249 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c249
*+ bl_0_249 br_0_249 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c249
*+ bl_0_249 br_0_249 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c249
*+ bl_0_249 br_0_249 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c249
*+ bl_0_249 br_0_249 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c249
*+ bl_0_249 br_0_249 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c249
*+ bl_0_249 br_0_249 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c249
*+ bl_0_249 br_0_249 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c249
*+ bl_0_249 br_0_249 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c249
*+ bl_0_249 br_0_249 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c249
*+ bl_0_249 br_0_249 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c249
*+ bl_0_249 br_0_249 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c249
*+ bl_0_249 br_0_249 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c249
*+ bl_0_249 br_0_249 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c249
*+ bl_0_249 br_0_249 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c249
*+ bl_0_249 br_0_249 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c249
*+ bl_0_249 br_0_249 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c249
*+ bl_0_249 br_0_249 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c249
*+ bl_0_249 br_0_249 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c249
*+ bl_0_249 br_0_249 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c249
*+ bl_0_249 br_0_249 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c249
*+ bl_0_249 br_0_249 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c249
*+ bl_0_249 br_0_249 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c249
*+ bl_0_249 br_0_249 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c249
*+ bl_0_249 br_0_249 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c249
*+ bl_0_249 br_0_249 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c249
*+ bl_0_249 br_0_249 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c249
*+ bl_0_249 br_0_249 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c249
*+ bl_0_249 br_0_249 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c249
*+ bl_0_249 br_0_249 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c249
*+ bl_0_249 br_0_249 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c249
*+ bl_0_249 br_0_249 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c249
*+ bl_0_249 br_0_249 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c249
*+ bl_0_249 br_0_249 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c249
*+ bl_0_249 br_0_249 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c249
*+ bl_0_249 br_0_249 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c249
*+ bl_0_249 br_0_249 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c249
*+ bl_0_249 br_0_249 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c249
*+ bl_0_249 br_0_249 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c249
*+ bl_0_249 br_0_249 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c249
*+ bl_0_249 br_0_249 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c249
*+ bl_0_249 br_0_249 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c249
*+ bl_0_249 br_0_249 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c249
*+ bl_0_249 br_0_249 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c249
*+ bl_0_249 br_0_249 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c249
*+ bl_0_249 br_0_249 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c249
*+ bl_0_249 br_0_249 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c249
*+ bl_0_249 br_0_249 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c249
*+ bl_0_249 br_0_249 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c249
*+ bl_0_249 br_0_249 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c249
*+ bl_0_249 br_0_249 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c249
*+ bl_0_249 br_0_249 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c249
*+ bl_0_249 br_0_249 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c249
*+ bl_0_249 br_0_249 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c249
*+ bl_0_249 br_0_249 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c249
*+ bl_0_249 br_0_249 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c249
*+ bl_0_249 br_0_249 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c249
*+ bl_0_249 br_0_249 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c249
*+ bl_0_249 br_0_249 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c249
*+ bl_0_249 br_0_249 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c249
*+ bl_0_249 br_0_249 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c249
*+ bl_0_249 br_0_249 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c249
*+ bl_0_249 br_0_249 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c249
*+ bl_0_249 br_0_249 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c249
*+ bl_0_249 br_0_249 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c249
*+ bl_0_249 br_0_249 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c249
*+ bl_0_249 br_0_249 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c249
*+ bl_0_249 br_0_249 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c249
*+ bl_0_249 br_0_249 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c249
*+ bl_0_249 br_0_249 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c249
*+ bl_0_249 br_0_249 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c249
*+ bl_0_249 br_0_249 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c249
*+ bl_0_249 br_0_249 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c249
*+ bl_0_249 br_0_249 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c249
*+ bl_0_249 br_0_249 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c249
*+ bl_0_249 br_0_249 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c249
*+ bl_0_249 br_0_249 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c249
*+ bl_0_249 br_0_249 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c249
*+ bl_0_249 br_0_249 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c249
+ bl_0_249 br_0_249 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c250
+ bl_0_250 br_0_250 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c250
*+ bl_0_250 br_0_250 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c250
*+ bl_0_250 br_0_250 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c250
*+ bl_0_250 br_0_250 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c250
*+ bl_0_250 br_0_250 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c250
*+ bl_0_250 br_0_250 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c250
*+ bl_0_250 br_0_250 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c250
*+ bl_0_250 br_0_250 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c250
*+ bl_0_250 br_0_250 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c250
*+ bl_0_250 br_0_250 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c250
*+ bl_0_250 br_0_250 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c250
*+ bl_0_250 br_0_250 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c250
*+ bl_0_250 br_0_250 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c250
*+ bl_0_250 br_0_250 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c250
*+ bl_0_250 br_0_250 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c250
*+ bl_0_250 br_0_250 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c250
*+ bl_0_250 br_0_250 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c250
*+ bl_0_250 br_0_250 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c250
*+ bl_0_250 br_0_250 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c250
*+ bl_0_250 br_0_250 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c250
*+ bl_0_250 br_0_250 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c250
*+ bl_0_250 br_0_250 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c250
*+ bl_0_250 br_0_250 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c250
*+ bl_0_250 br_0_250 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c250
*+ bl_0_250 br_0_250 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c250
*+ bl_0_250 br_0_250 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c250
*+ bl_0_250 br_0_250 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c250
*+ bl_0_250 br_0_250 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c250
*+ bl_0_250 br_0_250 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c250
*+ bl_0_250 br_0_250 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c250
*+ bl_0_250 br_0_250 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c250
*+ bl_0_250 br_0_250 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c250
*+ bl_0_250 br_0_250 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c250
*+ bl_0_250 br_0_250 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c250
*+ bl_0_250 br_0_250 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c250
*+ bl_0_250 br_0_250 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c250
*+ bl_0_250 br_0_250 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c250
*+ bl_0_250 br_0_250 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c250
*+ bl_0_250 br_0_250 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c250
*+ bl_0_250 br_0_250 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c250
*+ bl_0_250 br_0_250 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c250
*+ bl_0_250 br_0_250 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c250
*+ bl_0_250 br_0_250 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c250
*+ bl_0_250 br_0_250 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c250
*+ bl_0_250 br_0_250 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c250
*+ bl_0_250 br_0_250 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c250
*+ bl_0_250 br_0_250 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c250
*+ bl_0_250 br_0_250 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c250
*+ bl_0_250 br_0_250 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c250
*+ bl_0_250 br_0_250 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c250
*+ bl_0_250 br_0_250 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c250
*+ bl_0_250 br_0_250 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c250
*+ bl_0_250 br_0_250 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c250
*+ bl_0_250 br_0_250 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c250
*+ bl_0_250 br_0_250 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c250
*+ bl_0_250 br_0_250 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c250
*+ bl_0_250 br_0_250 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c250
*+ bl_0_250 br_0_250 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c250
*+ bl_0_250 br_0_250 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c250
*+ bl_0_250 br_0_250 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c250
*+ bl_0_250 br_0_250 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c250
*+ bl_0_250 br_0_250 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c250
*+ bl_0_250 br_0_250 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c250
*+ bl_0_250 br_0_250 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c250
*+ bl_0_250 br_0_250 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c250
*+ bl_0_250 br_0_250 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c250
*+ bl_0_250 br_0_250 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c250
*+ bl_0_250 br_0_250 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c250
*+ bl_0_250 br_0_250 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c250
*+ bl_0_250 br_0_250 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c250
*+ bl_0_250 br_0_250 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c250
*+ bl_0_250 br_0_250 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c250
*+ bl_0_250 br_0_250 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c250
*+ bl_0_250 br_0_250 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c250
*+ bl_0_250 br_0_250 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c250
*+ bl_0_250 br_0_250 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c250
*+ bl_0_250 br_0_250 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c250
*+ bl_0_250 br_0_250 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c250
*+ bl_0_250 br_0_250 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c250
*+ bl_0_250 br_0_250 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c250
*+ bl_0_250 br_0_250 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c250
*+ bl_0_250 br_0_250 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c250
*+ bl_0_250 br_0_250 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c250
*+ bl_0_250 br_0_250 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c250
*+ bl_0_250 br_0_250 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c250
*+ bl_0_250 br_0_250 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c250
*+ bl_0_250 br_0_250 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c250
*+ bl_0_250 br_0_250 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c250
*+ bl_0_250 br_0_250 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c250
*+ bl_0_250 br_0_250 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c250
*+ bl_0_250 br_0_250 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c250
*+ bl_0_250 br_0_250 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c250
*+ bl_0_250 br_0_250 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c250
*+ bl_0_250 br_0_250 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c250
*+ bl_0_250 br_0_250 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c250
*+ bl_0_250 br_0_250 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c250
*+ bl_0_250 br_0_250 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c250
*+ bl_0_250 br_0_250 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c250
*+ bl_0_250 br_0_250 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c250
*+ bl_0_250 br_0_250 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c250
*+ bl_0_250 br_0_250 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c250
*+ bl_0_250 br_0_250 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c250
*+ bl_0_250 br_0_250 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c250
*+ bl_0_250 br_0_250 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c250
*+ bl_0_250 br_0_250 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c250
*+ bl_0_250 br_0_250 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c250
*+ bl_0_250 br_0_250 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c250
*+ bl_0_250 br_0_250 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c250
*+ bl_0_250 br_0_250 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c250
*+ bl_0_250 br_0_250 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c250
*+ bl_0_250 br_0_250 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c250
*+ bl_0_250 br_0_250 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c250
*+ bl_0_250 br_0_250 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c250
*+ bl_0_250 br_0_250 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c250
*+ bl_0_250 br_0_250 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c250
*+ bl_0_250 br_0_250 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c250
*+ bl_0_250 br_0_250 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c250
*+ bl_0_250 br_0_250 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c250
*+ bl_0_250 br_0_250 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c250
*+ bl_0_250 br_0_250 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c250
*+ bl_0_250 br_0_250 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c250
*+ bl_0_250 br_0_250 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c250
*+ bl_0_250 br_0_250 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c250
*+ bl_0_250 br_0_250 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c250
*+ bl_0_250 br_0_250 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c250
*+ bl_0_250 br_0_250 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c250
*+ bl_0_250 br_0_250 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c250
+ bl_0_250 br_0_250 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c251
+ bl_0_251 br_0_251 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c251
*+ bl_0_251 br_0_251 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c251
*+ bl_0_251 br_0_251 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c251
*+ bl_0_251 br_0_251 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c251
*+ bl_0_251 br_0_251 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c251
*+ bl_0_251 br_0_251 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c251
*+ bl_0_251 br_0_251 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c251
*+ bl_0_251 br_0_251 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c251
*+ bl_0_251 br_0_251 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c251
*+ bl_0_251 br_0_251 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c251
*+ bl_0_251 br_0_251 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c251
*+ bl_0_251 br_0_251 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c251
*+ bl_0_251 br_0_251 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c251
*+ bl_0_251 br_0_251 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c251
*+ bl_0_251 br_0_251 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c251
*+ bl_0_251 br_0_251 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c251
*+ bl_0_251 br_0_251 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c251
*+ bl_0_251 br_0_251 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c251
*+ bl_0_251 br_0_251 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c251
*+ bl_0_251 br_0_251 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c251
*+ bl_0_251 br_0_251 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c251
*+ bl_0_251 br_0_251 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c251
*+ bl_0_251 br_0_251 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c251
*+ bl_0_251 br_0_251 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c251
*+ bl_0_251 br_0_251 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c251
*+ bl_0_251 br_0_251 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c251
*+ bl_0_251 br_0_251 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c251
*+ bl_0_251 br_0_251 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c251
*+ bl_0_251 br_0_251 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c251
*+ bl_0_251 br_0_251 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c251
*+ bl_0_251 br_0_251 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c251
*+ bl_0_251 br_0_251 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c251
*+ bl_0_251 br_0_251 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c251
*+ bl_0_251 br_0_251 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c251
*+ bl_0_251 br_0_251 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c251
*+ bl_0_251 br_0_251 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c251
*+ bl_0_251 br_0_251 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c251
*+ bl_0_251 br_0_251 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c251
*+ bl_0_251 br_0_251 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c251
*+ bl_0_251 br_0_251 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c251
*+ bl_0_251 br_0_251 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c251
*+ bl_0_251 br_0_251 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c251
*+ bl_0_251 br_0_251 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c251
*+ bl_0_251 br_0_251 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c251
*+ bl_0_251 br_0_251 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c251
*+ bl_0_251 br_0_251 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c251
*+ bl_0_251 br_0_251 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c251
*+ bl_0_251 br_0_251 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c251
*+ bl_0_251 br_0_251 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c251
*+ bl_0_251 br_0_251 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c251
*+ bl_0_251 br_0_251 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c251
*+ bl_0_251 br_0_251 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c251
*+ bl_0_251 br_0_251 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c251
*+ bl_0_251 br_0_251 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c251
*+ bl_0_251 br_0_251 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c251
*+ bl_0_251 br_0_251 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c251
*+ bl_0_251 br_0_251 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c251
*+ bl_0_251 br_0_251 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c251
*+ bl_0_251 br_0_251 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c251
*+ bl_0_251 br_0_251 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c251
*+ bl_0_251 br_0_251 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c251
*+ bl_0_251 br_0_251 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c251
*+ bl_0_251 br_0_251 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c251
*+ bl_0_251 br_0_251 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c251
*+ bl_0_251 br_0_251 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c251
*+ bl_0_251 br_0_251 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c251
*+ bl_0_251 br_0_251 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c251
*+ bl_0_251 br_0_251 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c251
*+ bl_0_251 br_0_251 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c251
*+ bl_0_251 br_0_251 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c251
*+ bl_0_251 br_0_251 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c251
*+ bl_0_251 br_0_251 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c251
*+ bl_0_251 br_0_251 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c251
*+ bl_0_251 br_0_251 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c251
*+ bl_0_251 br_0_251 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c251
*+ bl_0_251 br_0_251 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c251
*+ bl_0_251 br_0_251 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c251
*+ bl_0_251 br_0_251 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c251
*+ bl_0_251 br_0_251 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c251
*+ bl_0_251 br_0_251 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c251
*+ bl_0_251 br_0_251 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c251
*+ bl_0_251 br_0_251 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c251
*+ bl_0_251 br_0_251 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c251
*+ bl_0_251 br_0_251 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c251
*+ bl_0_251 br_0_251 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c251
*+ bl_0_251 br_0_251 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c251
*+ bl_0_251 br_0_251 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c251
*+ bl_0_251 br_0_251 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c251
*+ bl_0_251 br_0_251 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c251
*+ bl_0_251 br_0_251 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c251
*+ bl_0_251 br_0_251 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c251
*+ bl_0_251 br_0_251 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c251
*+ bl_0_251 br_0_251 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c251
*+ bl_0_251 br_0_251 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c251
*+ bl_0_251 br_0_251 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c251
*+ bl_0_251 br_0_251 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c251
*+ bl_0_251 br_0_251 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c251
*+ bl_0_251 br_0_251 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c251
*+ bl_0_251 br_0_251 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c251
*+ bl_0_251 br_0_251 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c251
*+ bl_0_251 br_0_251 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c251
*+ bl_0_251 br_0_251 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c251
*+ bl_0_251 br_0_251 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c251
*+ bl_0_251 br_0_251 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c251
*+ bl_0_251 br_0_251 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c251
*+ bl_0_251 br_0_251 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c251
*+ bl_0_251 br_0_251 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c251
*+ bl_0_251 br_0_251 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c251
*+ bl_0_251 br_0_251 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c251
*+ bl_0_251 br_0_251 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c251
*+ bl_0_251 br_0_251 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c251
*+ bl_0_251 br_0_251 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c251
*+ bl_0_251 br_0_251 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c251
*+ bl_0_251 br_0_251 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c251
*+ bl_0_251 br_0_251 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c251
*+ bl_0_251 br_0_251 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c251
*+ bl_0_251 br_0_251 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c251
*+ bl_0_251 br_0_251 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c251
*+ bl_0_251 br_0_251 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c251
*+ bl_0_251 br_0_251 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c251
*+ bl_0_251 br_0_251 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c251
*+ bl_0_251 br_0_251 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c251
*+ bl_0_251 br_0_251 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c251
*+ bl_0_251 br_0_251 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c251
*+ bl_0_251 br_0_251 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c251
*+ bl_0_251 br_0_251 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c251
*+ bl_0_251 br_0_251 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c251
+ bl_0_251 br_0_251 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c252
+ bl_0_252 br_0_252 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c252
*+ bl_0_252 br_0_252 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c252
*+ bl_0_252 br_0_252 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c252
*+ bl_0_252 br_0_252 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c252
*+ bl_0_252 br_0_252 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c252
*+ bl_0_252 br_0_252 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c252
*+ bl_0_252 br_0_252 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c252
*+ bl_0_252 br_0_252 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c252
*+ bl_0_252 br_0_252 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c252
*+ bl_0_252 br_0_252 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c252
*+ bl_0_252 br_0_252 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c252
*+ bl_0_252 br_0_252 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c252
*+ bl_0_252 br_0_252 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c252
*+ bl_0_252 br_0_252 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c252
*+ bl_0_252 br_0_252 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c252
*+ bl_0_252 br_0_252 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c252
*+ bl_0_252 br_0_252 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c252
*+ bl_0_252 br_0_252 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c252
*+ bl_0_252 br_0_252 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c252
*+ bl_0_252 br_0_252 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c252
*+ bl_0_252 br_0_252 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c252
*+ bl_0_252 br_0_252 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c252
*+ bl_0_252 br_0_252 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c252
*+ bl_0_252 br_0_252 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c252
*+ bl_0_252 br_0_252 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c252
*+ bl_0_252 br_0_252 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c252
*+ bl_0_252 br_0_252 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c252
*+ bl_0_252 br_0_252 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c252
*+ bl_0_252 br_0_252 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c252
*+ bl_0_252 br_0_252 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c252
*+ bl_0_252 br_0_252 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c252
*+ bl_0_252 br_0_252 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c252
*+ bl_0_252 br_0_252 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c252
*+ bl_0_252 br_0_252 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c252
*+ bl_0_252 br_0_252 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c252
*+ bl_0_252 br_0_252 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c252
*+ bl_0_252 br_0_252 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c252
*+ bl_0_252 br_0_252 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c252
*+ bl_0_252 br_0_252 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c252
*+ bl_0_252 br_0_252 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c252
*+ bl_0_252 br_0_252 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c252
*+ bl_0_252 br_0_252 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c252
*+ bl_0_252 br_0_252 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c252
*+ bl_0_252 br_0_252 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c252
*+ bl_0_252 br_0_252 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c252
*+ bl_0_252 br_0_252 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c252
*+ bl_0_252 br_0_252 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c252
*+ bl_0_252 br_0_252 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c252
*+ bl_0_252 br_0_252 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c252
*+ bl_0_252 br_0_252 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c252
*+ bl_0_252 br_0_252 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c252
*+ bl_0_252 br_0_252 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c252
*+ bl_0_252 br_0_252 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c252
*+ bl_0_252 br_0_252 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c252
*+ bl_0_252 br_0_252 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c252
*+ bl_0_252 br_0_252 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c252
*+ bl_0_252 br_0_252 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c252
*+ bl_0_252 br_0_252 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c252
*+ bl_0_252 br_0_252 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c252
*+ bl_0_252 br_0_252 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c252
*+ bl_0_252 br_0_252 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c252
*+ bl_0_252 br_0_252 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c252
*+ bl_0_252 br_0_252 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c252
*+ bl_0_252 br_0_252 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c252
*+ bl_0_252 br_0_252 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c252
*+ bl_0_252 br_0_252 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c252
*+ bl_0_252 br_0_252 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c252
*+ bl_0_252 br_0_252 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c252
*+ bl_0_252 br_0_252 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c252
*+ bl_0_252 br_0_252 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c252
*+ bl_0_252 br_0_252 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c252
*+ bl_0_252 br_0_252 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c252
*+ bl_0_252 br_0_252 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c252
*+ bl_0_252 br_0_252 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c252
*+ bl_0_252 br_0_252 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c252
*+ bl_0_252 br_0_252 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c252
*+ bl_0_252 br_0_252 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c252
*+ bl_0_252 br_0_252 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c252
*+ bl_0_252 br_0_252 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c252
*+ bl_0_252 br_0_252 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c252
*+ bl_0_252 br_0_252 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c252
*+ bl_0_252 br_0_252 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c252
*+ bl_0_252 br_0_252 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c252
*+ bl_0_252 br_0_252 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c252
*+ bl_0_252 br_0_252 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c252
*+ bl_0_252 br_0_252 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c252
*+ bl_0_252 br_0_252 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c252
*+ bl_0_252 br_0_252 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c252
*+ bl_0_252 br_0_252 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c252
*+ bl_0_252 br_0_252 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c252
*+ bl_0_252 br_0_252 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c252
*+ bl_0_252 br_0_252 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c252
*+ bl_0_252 br_0_252 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c252
*+ bl_0_252 br_0_252 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c252
*+ bl_0_252 br_0_252 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c252
*+ bl_0_252 br_0_252 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c252
*+ bl_0_252 br_0_252 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c252
*+ bl_0_252 br_0_252 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c252
*+ bl_0_252 br_0_252 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c252
*+ bl_0_252 br_0_252 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c252
*+ bl_0_252 br_0_252 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c252
*+ bl_0_252 br_0_252 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c252
*+ bl_0_252 br_0_252 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c252
*+ bl_0_252 br_0_252 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c252
*+ bl_0_252 br_0_252 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c252
*+ bl_0_252 br_0_252 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c252
*+ bl_0_252 br_0_252 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c252
*+ bl_0_252 br_0_252 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c252
*+ bl_0_252 br_0_252 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c252
*+ bl_0_252 br_0_252 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c252
*+ bl_0_252 br_0_252 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c252
*+ bl_0_252 br_0_252 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c252
*+ bl_0_252 br_0_252 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c252
*+ bl_0_252 br_0_252 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c252
*+ bl_0_252 br_0_252 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c252
*+ bl_0_252 br_0_252 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c252
*+ bl_0_252 br_0_252 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c252
*+ bl_0_252 br_0_252 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c252
*+ bl_0_252 br_0_252 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c252
*+ bl_0_252 br_0_252 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c252
*+ bl_0_252 br_0_252 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c252
*+ bl_0_252 br_0_252 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c252
*+ bl_0_252 br_0_252 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c252
*+ bl_0_252 br_0_252 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c252
*+ bl_0_252 br_0_252 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c252
*+ bl_0_252 br_0_252 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c252
*+ bl_0_252 br_0_252 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c252
+ bl_0_252 br_0_252 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c253
+ bl_0_253 br_0_253 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c253
*+ bl_0_253 br_0_253 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c253
*+ bl_0_253 br_0_253 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c253
*+ bl_0_253 br_0_253 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c253
*+ bl_0_253 br_0_253 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c253
*+ bl_0_253 br_0_253 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c253
*+ bl_0_253 br_0_253 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c253
*+ bl_0_253 br_0_253 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c253
*+ bl_0_253 br_0_253 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c253
*+ bl_0_253 br_0_253 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c253
*+ bl_0_253 br_0_253 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c253
*+ bl_0_253 br_0_253 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c253
*+ bl_0_253 br_0_253 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c253
*+ bl_0_253 br_0_253 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c253
*+ bl_0_253 br_0_253 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c253
*+ bl_0_253 br_0_253 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c253
*+ bl_0_253 br_0_253 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c253
*+ bl_0_253 br_0_253 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c253
*+ bl_0_253 br_0_253 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c253
*+ bl_0_253 br_0_253 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c253
*+ bl_0_253 br_0_253 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c253
*+ bl_0_253 br_0_253 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c253
*+ bl_0_253 br_0_253 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c253
*+ bl_0_253 br_0_253 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c253
*+ bl_0_253 br_0_253 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c253
*+ bl_0_253 br_0_253 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c253
*+ bl_0_253 br_0_253 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c253
*+ bl_0_253 br_0_253 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c253
*+ bl_0_253 br_0_253 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c253
*+ bl_0_253 br_0_253 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c253
*+ bl_0_253 br_0_253 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c253
*+ bl_0_253 br_0_253 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c253
*+ bl_0_253 br_0_253 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c253
*+ bl_0_253 br_0_253 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c253
*+ bl_0_253 br_0_253 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c253
*+ bl_0_253 br_0_253 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c253
*+ bl_0_253 br_0_253 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c253
*+ bl_0_253 br_0_253 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c253
*+ bl_0_253 br_0_253 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c253
*+ bl_0_253 br_0_253 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c253
*+ bl_0_253 br_0_253 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c253
*+ bl_0_253 br_0_253 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c253
*+ bl_0_253 br_0_253 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c253
*+ bl_0_253 br_0_253 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c253
*+ bl_0_253 br_0_253 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c253
*+ bl_0_253 br_0_253 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c253
*+ bl_0_253 br_0_253 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c253
*+ bl_0_253 br_0_253 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c253
*+ bl_0_253 br_0_253 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c253
*+ bl_0_253 br_0_253 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c253
*+ bl_0_253 br_0_253 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c253
*+ bl_0_253 br_0_253 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c253
*+ bl_0_253 br_0_253 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c253
*+ bl_0_253 br_0_253 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c253
*+ bl_0_253 br_0_253 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c253
*+ bl_0_253 br_0_253 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c253
*+ bl_0_253 br_0_253 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c253
*+ bl_0_253 br_0_253 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c253
*+ bl_0_253 br_0_253 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c253
*+ bl_0_253 br_0_253 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c253
*+ bl_0_253 br_0_253 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c253
*+ bl_0_253 br_0_253 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c253
*+ bl_0_253 br_0_253 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c253
*+ bl_0_253 br_0_253 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c253
*+ bl_0_253 br_0_253 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c253
*+ bl_0_253 br_0_253 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c253
*+ bl_0_253 br_0_253 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c253
*+ bl_0_253 br_0_253 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c253
*+ bl_0_253 br_0_253 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c253
*+ bl_0_253 br_0_253 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c253
*+ bl_0_253 br_0_253 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c253
*+ bl_0_253 br_0_253 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c253
*+ bl_0_253 br_0_253 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c253
*+ bl_0_253 br_0_253 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c253
*+ bl_0_253 br_0_253 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c253
*+ bl_0_253 br_0_253 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c253
*+ bl_0_253 br_0_253 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c253
*+ bl_0_253 br_0_253 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c253
*+ bl_0_253 br_0_253 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c253
*+ bl_0_253 br_0_253 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c253
*+ bl_0_253 br_0_253 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c253
*+ bl_0_253 br_0_253 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c253
*+ bl_0_253 br_0_253 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c253
*+ bl_0_253 br_0_253 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c253
*+ bl_0_253 br_0_253 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c253
*+ bl_0_253 br_0_253 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c253
*+ bl_0_253 br_0_253 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c253
*+ bl_0_253 br_0_253 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c253
*+ bl_0_253 br_0_253 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c253
*+ bl_0_253 br_0_253 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c253
*+ bl_0_253 br_0_253 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c253
*+ bl_0_253 br_0_253 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c253
*+ bl_0_253 br_0_253 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c253
*+ bl_0_253 br_0_253 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c253
*+ bl_0_253 br_0_253 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c253
*+ bl_0_253 br_0_253 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c253
*+ bl_0_253 br_0_253 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c253
*+ bl_0_253 br_0_253 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c253
*+ bl_0_253 br_0_253 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c253
*+ bl_0_253 br_0_253 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c253
*+ bl_0_253 br_0_253 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c253
*+ bl_0_253 br_0_253 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c253
*+ bl_0_253 br_0_253 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c253
*+ bl_0_253 br_0_253 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c253
*+ bl_0_253 br_0_253 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c253
*+ bl_0_253 br_0_253 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c253
*+ bl_0_253 br_0_253 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c253
*+ bl_0_253 br_0_253 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c253
*+ bl_0_253 br_0_253 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c253
*+ bl_0_253 br_0_253 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c253
*+ bl_0_253 br_0_253 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c253
*+ bl_0_253 br_0_253 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c253
*+ bl_0_253 br_0_253 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c253
*+ bl_0_253 br_0_253 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c253
*+ bl_0_253 br_0_253 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c253
*+ bl_0_253 br_0_253 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c253
*+ bl_0_253 br_0_253 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c253
*+ bl_0_253 br_0_253 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c253
*+ bl_0_253 br_0_253 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c253
*+ bl_0_253 br_0_253 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c253
*+ bl_0_253 br_0_253 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c253
*+ bl_0_253 br_0_253 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c253
*+ bl_0_253 br_0_253 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c253
*+ bl_0_253 br_0_253 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c253
*+ bl_0_253 br_0_253 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c253
*+ bl_0_253 br_0_253 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c253
*+ bl_0_253 br_0_253 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c253
+ bl_0_253 br_0_253 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c254
+ bl_0_254 br_0_254 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c254
*+ bl_0_254 br_0_254 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c254
*+ bl_0_254 br_0_254 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c254
*+ bl_0_254 br_0_254 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c254
*+ bl_0_254 br_0_254 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c254
*+ bl_0_254 br_0_254 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c254
*+ bl_0_254 br_0_254 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c254
*+ bl_0_254 br_0_254 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c254
*+ bl_0_254 br_0_254 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c254
*+ bl_0_254 br_0_254 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c254
*+ bl_0_254 br_0_254 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c254
*+ bl_0_254 br_0_254 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c254
*+ bl_0_254 br_0_254 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c254
*+ bl_0_254 br_0_254 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c254
*+ bl_0_254 br_0_254 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c254
*+ bl_0_254 br_0_254 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c254
*+ bl_0_254 br_0_254 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c254
*+ bl_0_254 br_0_254 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c254
*+ bl_0_254 br_0_254 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c254
*+ bl_0_254 br_0_254 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c254
*+ bl_0_254 br_0_254 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c254
*+ bl_0_254 br_0_254 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c254
*+ bl_0_254 br_0_254 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c254
*+ bl_0_254 br_0_254 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c254
*+ bl_0_254 br_0_254 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c254
*+ bl_0_254 br_0_254 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c254
*+ bl_0_254 br_0_254 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c254
*+ bl_0_254 br_0_254 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c254
*+ bl_0_254 br_0_254 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c254
*+ bl_0_254 br_0_254 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c254
*+ bl_0_254 br_0_254 wl_0_30 vdd gnd
*+ cell_1rw
* Xbit_r31_c254
*+ bl_0_254 br_0_254 wl_0_31 vdd gnd
*+ cell_1rw
* Xbit_r32_c254
*+ bl_0_254 br_0_254 wl_0_32 vdd gnd
*+ cell_1rw
* Xbit_r33_c254
*+ bl_0_254 br_0_254 wl_0_33 vdd gnd
*+ cell_1rw
* Xbit_r34_c254
*+ bl_0_254 br_0_254 wl_0_34 vdd gnd
*+ cell_1rw
* Xbit_r35_c254
*+ bl_0_254 br_0_254 wl_0_35 vdd gnd
*+ cell_1rw
* Xbit_r36_c254
*+ bl_0_254 br_0_254 wl_0_36 vdd gnd
*+ cell_1rw
* Xbit_r37_c254
*+ bl_0_254 br_0_254 wl_0_37 vdd gnd
*+ cell_1rw
* Xbit_r38_c254
*+ bl_0_254 br_0_254 wl_0_38 vdd gnd
*+ cell_1rw
* Xbit_r39_c254
*+ bl_0_254 br_0_254 wl_0_39 vdd gnd
*+ cell_1rw
* Xbit_r40_c254
*+ bl_0_254 br_0_254 wl_0_40 vdd gnd
*+ cell_1rw
* Xbit_r41_c254
*+ bl_0_254 br_0_254 wl_0_41 vdd gnd
*+ cell_1rw
* Xbit_r42_c254
*+ bl_0_254 br_0_254 wl_0_42 vdd gnd
*+ cell_1rw
* Xbit_r43_c254
*+ bl_0_254 br_0_254 wl_0_43 vdd gnd
*+ cell_1rw
* Xbit_r44_c254
*+ bl_0_254 br_0_254 wl_0_44 vdd gnd
*+ cell_1rw
* Xbit_r45_c254
*+ bl_0_254 br_0_254 wl_0_45 vdd gnd
*+ cell_1rw
* Xbit_r46_c254
*+ bl_0_254 br_0_254 wl_0_46 vdd gnd
*+ cell_1rw
* Xbit_r47_c254
*+ bl_0_254 br_0_254 wl_0_47 vdd gnd
*+ cell_1rw
* Xbit_r48_c254
*+ bl_0_254 br_0_254 wl_0_48 vdd gnd
*+ cell_1rw
* Xbit_r49_c254
*+ bl_0_254 br_0_254 wl_0_49 vdd gnd
*+ cell_1rw
* Xbit_r50_c254
*+ bl_0_254 br_0_254 wl_0_50 vdd gnd
*+ cell_1rw
* Xbit_r51_c254
*+ bl_0_254 br_0_254 wl_0_51 vdd gnd
*+ cell_1rw
* Xbit_r52_c254
*+ bl_0_254 br_0_254 wl_0_52 vdd gnd
*+ cell_1rw
* Xbit_r53_c254
*+ bl_0_254 br_0_254 wl_0_53 vdd gnd
*+ cell_1rw
* Xbit_r54_c254
*+ bl_0_254 br_0_254 wl_0_54 vdd gnd
*+ cell_1rw
* Xbit_r55_c254
*+ bl_0_254 br_0_254 wl_0_55 vdd gnd
*+ cell_1rw
* Xbit_r56_c254
*+ bl_0_254 br_0_254 wl_0_56 vdd gnd
*+ cell_1rw
* Xbit_r57_c254
*+ bl_0_254 br_0_254 wl_0_57 vdd gnd
*+ cell_1rw
* Xbit_r58_c254
*+ bl_0_254 br_0_254 wl_0_58 vdd gnd
*+ cell_1rw
* Xbit_r59_c254
*+ bl_0_254 br_0_254 wl_0_59 vdd gnd
*+ cell_1rw
* Xbit_r60_c254
*+ bl_0_254 br_0_254 wl_0_60 vdd gnd
*+ cell_1rw
* Xbit_r61_c254
*+ bl_0_254 br_0_254 wl_0_61 vdd gnd
*+ cell_1rw
* Xbit_r62_c254
*+ bl_0_254 br_0_254 wl_0_62 vdd gnd
*+ cell_1rw
* Xbit_r63_c254
*+ bl_0_254 br_0_254 wl_0_63 vdd gnd
*+ cell_1rw
* Xbit_r64_c254
*+ bl_0_254 br_0_254 wl_0_64 vdd gnd
*+ cell_1rw
* Xbit_r65_c254
*+ bl_0_254 br_0_254 wl_0_65 vdd gnd
*+ cell_1rw
* Xbit_r66_c254
*+ bl_0_254 br_0_254 wl_0_66 vdd gnd
*+ cell_1rw
* Xbit_r67_c254
*+ bl_0_254 br_0_254 wl_0_67 vdd gnd
*+ cell_1rw
* Xbit_r68_c254
*+ bl_0_254 br_0_254 wl_0_68 vdd gnd
*+ cell_1rw
* Xbit_r69_c254
*+ bl_0_254 br_0_254 wl_0_69 vdd gnd
*+ cell_1rw
* Xbit_r70_c254
*+ bl_0_254 br_0_254 wl_0_70 vdd gnd
*+ cell_1rw
* Xbit_r71_c254
*+ bl_0_254 br_0_254 wl_0_71 vdd gnd
*+ cell_1rw
* Xbit_r72_c254
*+ bl_0_254 br_0_254 wl_0_72 vdd gnd
*+ cell_1rw
* Xbit_r73_c254
*+ bl_0_254 br_0_254 wl_0_73 vdd gnd
*+ cell_1rw
* Xbit_r74_c254
*+ bl_0_254 br_0_254 wl_0_74 vdd gnd
*+ cell_1rw
* Xbit_r75_c254
*+ bl_0_254 br_0_254 wl_0_75 vdd gnd
*+ cell_1rw
* Xbit_r76_c254
*+ bl_0_254 br_0_254 wl_0_76 vdd gnd
*+ cell_1rw
* Xbit_r77_c254
*+ bl_0_254 br_0_254 wl_0_77 vdd gnd
*+ cell_1rw
* Xbit_r78_c254
*+ bl_0_254 br_0_254 wl_0_78 vdd gnd
*+ cell_1rw
* Xbit_r79_c254
*+ bl_0_254 br_0_254 wl_0_79 vdd gnd
*+ cell_1rw
* Xbit_r80_c254
*+ bl_0_254 br_0_254 wl_0_80 vdd gnd
*+ cell_1rw
* Xbit_r81_c254
*+ bl_0_254 br_0_254 wl_0_81 vdd gnd
*+ cell_1rw
* Xbit_r82_c254
*+ bl_0_254 br_0_254 wl_0_82 vdd gnd
*+ cell_1rw
* Xbit_r83_c254
*+ bl_0_254 br_0_254 wl_0_83 vdd gnd
*+ cell_1rw
* Xbit_r84_c254
*+ bl_0_254 br_0_254 wl_0_84 vdd gnd
*+ cell_1rw
* Xbit_r85_c254
*+ bl_0_254 br_0_254 wl_0_85 vdd gnd
*+ cell_1rw
* Xbit_r86_c254
*+ bl_0_254 br_0_254 wl_0_86 vdd gnd
*+ cell_1rw
* Xbit_r87_c254
*+ bl_0_254 br_0_254 wl_0_87 vdd gnd
*+ cell_1rw
* Xbit_r88_c254
*+ bl_0_254 br_0_254 wl_0_88 vdd gnd
*+ cell_1rw
* Xbit_r89_c254
*+ bl_0_254 br_0_254 wl_0_89 vdd gnd
*+ cell_1rw
* Xbit_r90_c254
*+ bl_0_254 br_0_254 wl_0_90 vdd gnd
*+ cell_1rw
* Xbit_r91_c254
*+ bl_0_254 br_0_254 wl_0_91 vdd gnd
*+ cell_1rw
* Xbit_r92_c254
*+ bl_0_254 br_0_254 wl_0_92 vdd gnd
*+ cell_1rw
* Xbit_r93_c254
*+ bl_0_254 br_0_254 wl_0_93 vdd gnd
*+ cell_1rw
* Xbit_r94_c254
*+ bl_0_254 br_0_254 wl_0_94 vdd gnd
*+ cell_1rw
* Xbit_r95_c254
*+ bl_0_254 br_0_254 wl_0_95 vdd gnd
*+ cell_1rw
* Xbit_r96_c254
*+ bl_0_254 br_0_254 wl_0_96 vdd gnd
*+ cell_1rw
* Xbit_r97_c254
*+ bl_0_254 br_0_254 wl_0_97 vdd gnd
*+ cell_1rw
* Xbit_r98_c254
*+ bl_0_254 br_0_254 wl_0_98 vdd gnd
*+ cell_1rw
* Xbit_r99_c254
*+ bl_0_254 br_0_254 wl_0_99 vdd gnd
*+ cell_1rw
* Xbit_r100_c254
*+ bl_0_254 br_0_254 wl_0_100 vdd gnd
*+ cell_1rw
* Xbit_r101_c254
*+ bl_0_254 br_0_254 wl_0_101 vdd gnd
*+ cell_1rw
* Xbit_r102_c254
*+ bl_0_254 br_0_254 wl_0_102 vdd gnd
*+ cell_1rw
* Xbit_r103_c254
*+ bl_0_254 br_0_254 wl_0_103 vdd gnd
*+ cell_1rw
* Xbit_r104_c254
*+ bl_0_254 br_0_254 wl_0_104 vdd gnd
*+ cell_1rw
* Xbit_r105_c254
*+ bl_0_254 br_0_254 wl_0_105 vdd gnd
*+ cell_1rw
* Xbit_r106_c254
*+ bl_0_254 br_0_254 wl_0_106 vdd gnd
*+ cell_1rw
* Xbit_r107_c254
*+ bl_0_254 br_0_254 wl_0_107 vdd gnd
*+ cell_1rw
* Xbit_r108_c254
*+ bl_0_254 br_0_254 wl_0_108 vdd gnd
*+ cell_1rw
* Xbit_r109_c254
*+ bl_0_254 br_0_254 wl_0_109 vdd gnd
*+ cell_1rw
* Xbit_r110_c254
*+ bl_0_254 br_0_254 wl_0_110 vdd gnd
*+ cell_1rw
* Xbit_r111_c254
*+ bl_0_254 br_0_254 wl_0_111 vdd gnd
*+ cell_1rw
* Xbit_r112_c254
*+ bl_0_254 br_0_254 wl_0_112 vdd gnd
*+ cell_1rw
* Xbit_r113_c254
*+ bl_0_254 br_0_254 wl_0_113 vdd gnd
*+ cell_1rw
* Xbit_r114_c254
*+ bl_0_254 br_0_254 wl_0_114 vdd gnd
*+ cell_1rw
* Xbit_r115_c254
*+ bl_0_254 br_0_254 wl_0_115 vdd gnd
*+ cell_1rw
* Xbit_r116_c254
*+ bl_0_254 br_0_254 wl_0_116 vdd gnd
*+ cell_1rw
* Xbit_r117_c254
*+ bl_0_254 br_0_254 wl_0_117 vdd gnd
*+ cell_1rw
* Xbit_r118_c254
*+ bl_0_254 br_0_254 wl_0_118 vdd gnd
*+ cell_1rw
* Xbit_r119_c254
*+ bl_0_254 br_0_254 wl_0_119 vdd gnd
*+ cell_1rw
* Xbit_r120_c254
*+ bl_0_254 br_0_254 wl_0_120 vdd gnd
*+ cell_1rw
* Xbit_r121_c254
*+ bl_0_254 br_0_254 wl_0_121 vdd gnd
*+ cell_1rw
* Xbit_r122_c254
*+ bl_0_254 br_0_254 wl_0_122 vdd gnd
*+ cell_1rw
* Xbit_r123_c254
*+ bl_0_254 br_0_254 wl_0_123 vdd gnd
*+ cell_1rw
* Xbit_r124_c254
*+ bl_0_254 br_0_254 wl_0_124 vdd gnd
*+ cell_1rw
* Xbit_r125_c254
*+ bl_0_254 br_0_254 wl_0_125 vdd gnd
*+ cell_1rw
* Xbit_r126_c254
*+ bl_0_254 br_0_254 wl_0_126 vdd gnd
*+ cell_1rw
Xbit_r127_c254
+ bl_0_254 br_0_254 wl_0_127 vdd gnd
+ cell_1rw
Xbit_r0_c255
+ bl_0_255 br_0_255 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c255
+ bl_0_255 br_0_255 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c255
+ bl_0_255 br_0_255 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c255
+ bl_0_255 br_0_255 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c255
+ bl_0_255 br_0_255 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c255
+ bl_0_255 br_0_255 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c255
+ bl_0_255 br_0_255 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c255
+ bl_0_255 br_0_255 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c255
+ bl_0_255 br_0_255 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c255
+ bl_0_255 br_0_255 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c255
+ bl_0_255 br_0_255 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c255
+ bl_0_255 br_0_255 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c255
+ bl_0_255 br_0_255 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c255
+ bl_0_255 br_0_255 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c255
+ bl_0_255 br_0_255 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c255
+ bl_0_255 br_0_255 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c255
+ bl_0_255 br_0_255 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c255
+ bl_0_255 br_0_255 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c255
+ bl_0_255 br_0_255 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c255
+ bl_0_255 br_0_255 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c255
+ bl_0_255 br_0_255 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c255
+ bl_0_255 br_0_255 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c255
+ bl_0_255 br_0_255 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c255
+ bl_0_255 br_0_255 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c255
+ bl_0_255 br_0_255 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c255
+ bl_0_255 br_0_255 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c255
+ bl_0_255 br_0_255 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c255
+ bl_0_255 br_0_255 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c255
+ bl_0_255 br_0_255 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c255
+ bl_0_255 br_0_255 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c255
+ bl_0_255 br_0_255 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c255
+ bl_0_255 br_0_255 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r32_c255
+ bl_0_255 br_0_255 wl_0_32 vdd gnd
+ cell_1rw
Xbit_r33_c255
+ bl_0_255 br_0_255 wl_0_33 vdd gnd
+ cell_1rw
Xbit_r34_c255
+ bl_0_255 br_0_255 wl_0_34 vdd gnd
+ cell_1rw
Xbit_r35_c255
+ bl_0_255 br_0_255 wl_0_35 vdd gnd
+ cell_1rw
Xbit_r36_c255
+ bl_0_255 br_0_255 wl_0_36 vdd gnd
+ cell_1rw
Xbit_r37_c255
+ bl_0_255 br_0_255 wl_0_37 vdd gnd
+ cell_1rw
Xbit_r38_c255
+ bl_0_255 br_0_255 wl_0_38 vdd gnd
+ cell_1rw
Xbit_r39_c255
+ bl_0_255 br_0_255 wl_0_39 vdd gnd
+ cell_1rw
Xbit_r40_c255
+ bl_0_255 br_0_255 wl_0_40 vdd gnd
+ cell_1rw
Xbit_r41_c255
+ bl_0_255 br_0_255 wl_0_41 vdd gnd
+ cell_1rw
Xbit_r42_c255
+ bl_0_255 br_0_255 wl_0_42 vdd gnd
+ cell_1rw
Xbit_r43_c255
+ bl_0_255 br_0_255 wl_0_43 vdd gnd
+ cell_1rw
Xbit_r44_c255
+ bl_0_255 br_0_255 wl_0_44 vdd gnd
+ cell_1rw
Xbit_r45_c255
+ bl_0_255 br_0_255 wl_0_45 vdd gnd
+ cell_1rw
Xbit_r46_c255
+ bl_0_255 br_0_255 wl_0_46 vdd gnd
+ cell_1rw
Xbit_r47_c255
+ bl_0_255 br_0_255 wl_0_47 vdd gnd
+ cell_1rw
Xbit_r48_c255
+ bl_0_255 br_0_255 wl_0_48 vdd gnd
+ cell_1rw
Xbit_r49_c255
+ bl_0_255 br_0_255 wl_0_49 vdd gnd
+ cell_1rw
Xbit_r50_c255
+ bl_0_255 br_0_255 wl_0_50 vdd gnd
+ cell_1rw
Xbit_r51_c255
+ bl_0_255 br_0_255 wl_0_51 vdd gnd
+ cell_1rw
Xbit_r52_c255
+ bl_0_255 br_0_255 wl_0_52 vdd gnd
+ cell_1rw
Xbit_r53_c255
+ bl_0_255 br_0_255 wl_0_53 vdd gnd
+ cell_1rw
Xbit_r54_c255
+ bl_0_255 br_0_255 wl_0_54 vdd gnd
+ cell_1rw
Xbit_r55_c255
+ bl_0_255 br_0_255 wl_0_55 vdd gnd
+ cell_1rw
Xbit_r56_c255
+ bl_0_255 br_0_255 wl_0_56 vdd gnd
+ cell_1rw
Xbit_r57_c255
+ bl_0_255 br_0_255 wl_0_57 vdd gnd
+ cell_1rw
Xbit_r58_c255
+ bl_0_255 br_0_255 wl_0_58 vdd gnd
+ cell_1rw
Xbit_r59_c255
+ bl_0_255 br_0_255 wl_0_59 vdd gnd
+ cell_1rw
Xbit_r60_c255
+ bl_0_255 br_0_255 wl_0_60 vdd gnd
+ cell_1rw
Xbit_r61_c255
+ bl_0_255 br_0_255 wl_0_61 vdd gnd
+ cell_1rw
Xbit_r62_c255
+ bl_0_255 br_0_255 wl_0_62 vdd gnd
+ cell_1rw
Xbit_r63_c255
+ bl_0_255 br_0_255 wl_0_63 vdd gnd
+ cell_1rw
Xbit_r64_c255
+ bl_0_255 br_0_255 wl_0_64 vdd gnd
+ cell_1rw
Xbit_r65_c255
+ bl_0_255 br_0_255 wl_0_65 vdd gnd
+ cell_1rw
Xbit_r66_c255
+ bl_0_255 br_0_255 wl_0_66 vdd gnd
+ cell_1rw
Xbit_r67_c255
+ bl_0_255 br_0_255 wl_0_67 vdd gnd
+ cell_1rw
Xbit_r68_c255
+ bl_0_255 br_0_255 wl_0_68 vdd gnd
+ cell_1rw
Xbit_r69_c255
+ bl_0_255 br_0_255 wl_0_69 vdd gnd
+ cell_1rw
Xbit_r70_c255
+ bl_0_255 br_0_255 wl_0_70 vdd gnd
+ cell_1rw
Xbit_r71_c255
+ bl_0_255 br_0_255 wl_0_71 vdd gnd
+ cell_1rw
Xbit_r72_c255
+ bl_0_255 br_0_255 wl_0_72 vdd gnd
+ cell_1rw
Xbit_r73_c255
+ bl_0_255 br_0_255 wl_0_73 vdd gnd
+ cell_1rw
Xbit_r74_c255
+ bl_0_255 br_0_255 wl_0_74 vdd gnd
+ cell_1rw
Xbit_r75_c255
+ bl_0_255 br_0_255 wl_0_75 vdd gnd
+ cell_1rw
Xbit_r76_c255
+ bl_0_255 br_0_255 wl_0_76 vdd gnd
+ cell_1rw
Xbit_r77_c255
+ bl_0_255 br_0_255 wl_0_77 vdd gnd
+ cell_1rw
Xbit_r78_c255
+ bl_0_255 br_0_255 wl_0_78 vdd gnd
+ cell_1rw
Xbit_r79_c255
+ bl_0_255 br_0_255 wl_0_79 vdd gnd
+ cell_1rw
Xbit_r80_c255
+ bl_0_255 br_0_255 wl_0_80 vdd gnd
+ cell_1rw
Xbit_r81_c255
+ bl_0_255 br_0_255 wl_0_81 vdd gnd
+ cell_1rw
Xbit_r82_c255
+ bl_0_255 br_0_255 wl_0_82 vdd gnd
+ cell_1rw
Xbit_r83_c255
+ bl_0_255 br_0_255 wl_0_83 vdd gnd
+ cell_1rw
Xbit_r84_c255
+ bl_0_255 br_0_255 wl_0_84 vdd gnd
+ cell_1rw
Xbit_r85_c255
+ bl_0_255 br_0_255 wl_0_85 vdd gnd
+ cell_1rw
Xbit_r86_c255
+ bl_0_255 br_0_255 wl_0_86 vdd gnd
+ cell_1rw
Xbit_r87_c255
+ bl_0_255 br_0_255 wl_0_87 vdd gnd
+ cell_1rw
Xbit_r88_c255
+ bl_0_255 br_0_255 wl_0_88 vdd gnd
+ cell_1rw
Xbit_r89_c255
+ bl_0_255 br_0_255 wl_0_89 vdd gnd
+ cell_1rw
Xbit_r90_c255
+ bl_0_255 br_0_255 wl_0_90 vdd gnd
+ cell_1rw
Xbit_r91_c255
+ bl_0_255 br_0_255 wl_0_91 vdd gnd
+ cell_1rw
Xbit_r92_c255
+ bl_0_255 br_0_255 wl_0_92 vdd gnd
+ cell_1rw
Xbit_r93_c255
+ bl_0_255 br_0_255 wl_0_93 vdd gnd
+ cell_1rw
Xbit_r94_c255
+ bl_0_255 br_0_255 wl_0_94 vdd gnd
+ cell_1rw
Xbit_r95_c255
+ bl_0_255 br_0_255 wl_0_95 vdd gnd
+ cell_1rw
Xbit_r96_c255
+ bl_0_255 br_0_255 wl_0_96 vdd gnd
+ cell_1rw
Xbit_r97_c255
+ bl_0_255 br_0_255 wl_0_97 vdd gnd
+ cell_1rw
Xbit_r98_c255
+ bl_0_255 br_0_255 wl_0_98 vdd gnd
+ cell_1rw
Xbit_r99_c255
+ bl_0_255 br_0_255 wl_0_99 vdd gnd
+ cell_1rw
Xbit_r100_c255
+ bl_0_255 br_0_255 wl_0_100 vdd gnd
+ cell_1rw
Xbit_r101_c255
+ bl_0_255 br_0_255 wl_0_101 vdd gnd
+ cell_1rw
Xbit_r102_c255
+ bl_0_255 br_0_255 wl_0_102 vdd gnd
+ cell_1rw
Xbit_r103_c255
+ bl_0_255 br_0_255 wl_0_103 vdd gnd
+ cell_1rw
Xbit_r104_c255
+ bl_0_255 br_0_255 wl_0_104 vdd gnd
+ cell_1rw
Xbit_r105_c255
+ bl_0_255 br_0_255 wl_0_105 vdd gnd
+ cell_1rw
Xbit_r106_c255
+ bl_0_255 br_0_255 wl_0_106 vdd gnd
+ cell_1rw
Xbit_r107_c255
+ bl_0_255 br_0_255 wl_0_107 vdd gnd
+ cell_1rw
Xbit_r108_c255
+ bl_0_255 br_0_255 wl_0_108 vdd gnd
+ cell_1rw
Xbit_r109_c255
+ bl_0_255 br_0_255 wl_0_109 vdd gnd
+ cell_1rw
Xbit_r110_c255
+ bl_0_255 br_0_255 wl_0_110 vdd gnd
+ cell_1rw
Xbit_r111_c255
+ bl_0_255 br_0_255 wl_0_111 vdd gnd
+ cell_1rw
Xbit_r112_c255
+ bl_0_255 br_0_255 wl_0_112 vdd gnd
+ cell_1rw
Xbit_r113_c255
+ bl_0_255 br_0_255 wl_0_113 vdd gnd
+ cell_1rw
Xbit_r114_c255
+ bl_0_255 br_0_255 wl_0_114 vdd gnd
+ cell_1rw
Xbit_r115_c255
+ bl_0_255 br_0_255 wl_0_115 vdd gnd
+ cell_1rw
Xbit_r116_c255
+ bl_0_255 br_0_255 wl_0_116 vdd gnd
+ cell_1rw
Xbit_r117_c255
+ bl_0_255 br_0_255 wl_0_117 vdd gnd
+ cell_1rw
Xbit_r118_c255
+ bl_0_255 br_0_255 wl_0_118 vdd gnd
+ cell_1rw
Xbit_r119_c255
+ bl_0_255 br_0_255 wl_0_119 vdd gnd
+ cell_1rw
Xbit_r120_c255
+ bl_0_255 br_0_255 wl_0_120 vdd gnd
+ cell_1rw
Xbit_r121_c255
+ bl_0_255 br_0_255 wl_0_121 vdd gnd
+ cell_1rw
Xbit_r122_c255
+ bl_0_255 br_0_255 wl_0_122 vdd gnd
+ cell_1rw
Xbit_r123_c255
+ bl_0_255 br_0_255 wl_0_123 vdd gnd
+ cell_1rw
Xbit_r124_c255
+ bl_0_255 br_0_255 wl_0_124 vdd gnd
+ cell_1rw
Xbit_r125_c255
+ bl_0_255 br_0_255 wl_0_125 vdd gnd
+ cell_1rw
Xbit_r126_c255
+ bl_0_255 br_0_255 wl_0_126 vdd gnd
+ cell_1rw
Xbit_r127_c255
+ bl_0_255 br_0_255 wl_0_127 vdd gnd
+ cell_1rw
.ENDS sram_1rw0r0w_32_1024_freepdk45_bitcell_array

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_replica_bitcell_array
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64
+ bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68
+ bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72
+ bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76
+ bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80
+ bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84
+ bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88
+ bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92
+ bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96
+ bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100
+ bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104
+ br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107
+ bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111
+ br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114
+ bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118
+ br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121
+ bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125
+ br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128
+ bl_0_129 br_0_129 bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132
+ br_0_132 bl_0_133 br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135
+ bl_0_136 br_0_136 bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139
+ br_0_139 bl_0_140 br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142
+ bl_0_143 br_0_143 bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146
+ br_0_146 bl_0_147 br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149
+ bl_0_150 br_0_150 bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153
+ br_0_153 bl_0_154 br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156
+ bl_0_157 br_0_157 bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160
+ br_0_160 bl_0_161 br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163
+ bl_0_164 br_0_164 bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167
+ br_0_167 bl_0_168 br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170
+ bl_0_171 br_0_171 bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174
+ br_0_174 bl_0_175 br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177
+ bl_0_178 br_0_178 bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181
+ br_0_181 bl_0_182 br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184
+ bl_0_185 br_0_185 bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188
+ br_0_188 bl_0_189 br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191
+ bl_0_192 br_0_192 bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195
+ br_0_195 bl_0_196 br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198
+ bl_0_199 br_0_199 bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202
+ br_0_202 bl_0_203 br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205
+ bl_0_206 br_0_206 bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209
+ br_0_209 bl_0_210 br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212
+ bl_0_213 br_0_213 bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216
+ br_0_216 bl_0_217 br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219
+ bl_0_220 br_0_220 bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223
+ br_0_223 bl_0_224 br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226
+ bl_0_227 br_0_227 bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230
+ br_0_230 bl_0_231 br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233
+ bl_0_234 br_0_234 bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237
+ br_0_237 bl_0_238 br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240
+ bl_0_241 br_0_241 bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244
+ br_0_244 bl_0_245 br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247
+ bl_0_248 br_0_248 bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251
+ br_0_251 bl_0_252 br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254
+ bl_0_255 br_0_255 rbl_wl_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5
+ wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14
+ wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22
+ wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30
+ wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38
+ wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46
+ wl_0_47 wl_0_48 wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54
+ wl_0_55 wl_0_56 wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62
+ wl_0_63 wl_0_64 wl_0_65 wl_0_66 wl_0_67 wl_0_68 wl_0_69 wl_0_70
+ wl_0_71 wl_0_72 wl_0_73 wl_0_74 wl_0_75 wl_0_76 wl_0_77 wl_0_78
+ wl_0_79 wl_0_80 wl_0_81 wl_0_82 wl_0_83 wl_0_84 wl_0_85 wl_0_86
+ wl_0_87 wl_0_88 wl_0_89 wl_0_90 wl_0_91 wl_0_92 wl_0_93 wl_0_94
+ wl_0_95 wl_0_96 wl_0_97 wl_0_98 wl_0_99 wl_0_100 wl_0_101 wl_0_102
+ wl_0_103 wl_0_104 wl_0_105 wl_0_106 wl_0_107 wl_0_108 wl_0_109
+ wl_0_110 wl_0_111 wl_0_112 wl_0_113 wl_0_114 wl_0_115 wl_0_116
+ wl_0_117 wl_0_118 wl_0_119 wl_0_120 wl_0_121 wl_0_122 wl_0_123
+ wl_0_124 wl_0_125 wl_0_126 wl_0_127 vdd gnd
* INOUT : rbl_bl_0_0 
* INOUT : rbl_br_0_0 
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INOUT : bl_0_64 
* INOUT : br_0_64 
* INOUT : bl_0_65 
* INOUT : br_0_65 
* INOUT : bl_0_66 
* INOUT : br_0_66 
* INOUT : bl_0_67 
* INOUT : br_0_67 
* INOUT : bl_0_68 
* INOUT : br_0_68 
* INOUT : bl_0_69 
* INOUT : br_0_69 
* INOUT : bl_0_70 
* INOUT : br_0_70 
* INOUT : bl_0_71 
* INOUT : br_0_71 
* INOUT : bl_0_72 
* INOUT : br_0_72 
* INOUT : bl_0_73 
* INOUT : br_0_73 
* INOUT : bl_0_74 
* INOUT : br_0_74 
* INOUT : bl_0_75 
* INOUT : br_0_75 
* INOUT : bl_0_76 
* INOUT : br_0_76 
* INOUT : bl_0_77 
* INOUT : br_0_77 
* INOUT : bl_0_78 
* INOUT : br_0_78 
* INOUT : bl_0_79 
* INOUT : br_0_79 
* INOUT : bl_0_80 
* INOUT : br_0_80 
* INOUT : bl_0_81 
* INOUT : br_0_81 
* INOUT : bl_0_82 
* INOUT : br_0_82 
* INOUT : bl_0_83 
* INOUT : br_0_83 
* INOUT : bl_0_84 
* INOUT : br_0_84 
* INOUT : bl_0_85 
* INOUT : br_0_85 
* INOUT : bl_0_86 
* INOUT : br_0_86 
* INOUT : bl_0_87 
* INOUT : br_0_87 
* INOUT : bl_0_88 
* INOUT : br_0_88 
* INOUT : bl_0_89 
* INOUT : br_0_89 
* INOUT : bl_0_90 
* INOUT : br_0_90 
* INOUT : bl_0_91 
* INOUT : br_0_91 
* INOUT : bl_0_92 
* INOUT : br_0_92 
* INOUT : bl_0_93 
* INOUT : br_0_93 
* INOUT : bl_0_94 
* INOUT : br_0_94 
* INOUT : bl_0_95 
* INOUT : br_0_95 
* INOUT : bl_0_96 
* INOUT : br_0_96 
* INOUT : bl_0_97 
* INOUT : br_0_97 
* INOUT : bl_0_98 
* INOUT : br_0_98 
* INOUT : bl_0_99 
* INOUT : br_0_99 
* INOUT : bl_0_100 
* INOUT : br_0_100 
* INOUT : bl_0_101 
* INOUT : br_0_101 
* INOUT : bl_0_102 
* INOUT : br_0_102 
* INOUT : bl_0_103 
* INOUT : br_0_103 
* INOUT : bl_0_104 
* INOUT : br_0_104 
* INOUT : bl_0_105 
* INOUT : br_0_105 
* INOUT : bl_0_106 
* INOUT : br_0_106 
* INOUT : bl_0_107 
* INOUT : br_0_107 
* INOUT : bl_0_108 
* INOUT : br_0_108 
* INOUT : bl_0_109 
* INOUT : br_0_109 
* INOUT : bl_0_110 
* INOUT : br_0_110 
* INOUT : bl_0_111 
* INOUT : br_0_111 
* INOUT : bl_0_112 
* INOUT : br_0_112 
* INOUT : bl_0_113 
* INOUT : br_0_113 
* INOUT : bl_0_114 
* INOUT : br_0_114 
* INOUT : bl_0_115 
* INOUT : br_0_115 
* INOUT : bl_0_116 
* INOUT : br_0_116 
* INOUT : bl_0_117 
* INOUT : br_0_117 
* INOUT : bl_0_118 
* INOUT : br_0_118 
* INOUT : bl_0_119 
* INOUT : br_0_119 
* INOUT : bl_0_120 
* INOUT : br_0_120 
* INOUT : bl_0_121 
* INOUT : br_0_121 
* INOUT : bl_0_122 
* INOUT : br_0_122 
* INOUT : bl_0_123 
* INOUT : br_0_123 
* INOUT : bl_0_124 
* INOUT : br_0_124 
* INOUT : bl_0_125 
* INOUT : br_0_125 
* INOUT : bl_0_126 
* INOUT : br_0_126 
* INOUT : bl_0_127 
* INOUT : br_0_127 
* INOUT : bl_0_128 
* INOUT : br_0_128 
* INOUT : bl_0_129 
* INOUT : br_0_129 
* INOUT : bl_0_130 
* INOUT : br_0_130 
* INOUT : bl_0_131 
* INOUT : br_0_131 
* INOUT : bl_0_132 
* INOUT : br_0_132 
* INOUT : bl_0_133 
* INOUT : br_0_133 
* INOUT : bl_0_134 
* INOUT : br_0_134 
* INOUT : bl_0_135 
* INOUT : br_0_135 
* INOUT : bl_0_136 
* INOUT : br_0_136 
* INOUT : bl_0_137 
* INOUT : br_0_137 
* INOUT : bl_0_138 
* INOUT : br_0_138 
* INOUT : bl_0_139 
* INOUT : br_0_139 
* INOUT : bl_0_140 
* INOUT : br_0_140 
* INOUT : bl_0_141 
* INOUT : br_0_141 
* INOUT : bl_0_142 
* INOUT : br_0_142 
* INOUT : bl_0_143 
* INOUT : br_0_143 
* INOUT : bl_0_144 
* INOUT : br_0_144 
* INOUT : bl_0_145 
* INOUT : br_0_145 
* INOUT : bl_0_146 
* INOUT : br_0_146 
* INOUT : bl_0_147 
* INOUT : br_0_147 
* INOUT : bl_0_148 
* INOUT : br_0_148 
* INOUT : bl_0_149 
* INOUT : br_0_149 
* INOUT : bl_0_150 
* INOUT : br_0_150 
* INOUT : bl_0_151 
* INOUT : br_0_151 
* INOUT : bl_0_152 
* INOUT : br_0_152 
* INOUT : bl_0_153 
* INOUT : br_0_153 
* INOUT : bl_0_154 
* INOUT : br_0_154 
* INOUT : bl_0_155 
* INOUT : br_0_155 
* INOUT : bl_0_156 
* INOUT : br_0_156 
* INOUT : bl_0_157 
* INOUT : br_0_157 
* INOUT : bl_0_158 
* INOUT : br_0_158 
* INOUT : bl_0_159 
* INOUT : br_0_159 
* INOUT : bl_0_160 
* INOUT : br_0_160 
* INOUT : bl_0_161 
* INOUT : br_0_161 
* INOUT : bl_0_162 
* INOUT : br_0_162 
* INOUT : bl_0_163 
* INOUT : br_0_163 
* INOUT : bl_0_164 
* INOUT : br_0_164 
* INOUT : bl_0_165 
* INOUT : br_0_165 
* INOUT : bl_0_166 
* INOUT : br_0_166 
* INOUT : bl_0_167 
* INOUT : br_0_167 
* INOUT : bl_0_168 
* INOUT : br_0_168 
* INOUT : bl_0_169 
* INOUT : br_0_169 
* INOUT : bl_0_170 
* INOUT : br_0_170 
* INOUT : bl_0_171 
* INOUT : br_0_171 
* INOUT : bl_0_172 
* INOUT : br_0_172 
* INOUT : bl_0_173 
* INOUT : br_0_173 
* INOUT : bl_0_174 
* INOUT : br_0_174 
* INOUT : bl_0_175 
* INOUT : br_0_175 
* INOUT : bl_0_176 
* INOUT : br_0_176 
* INOUT : bl_0_177 
* INOUT : br_0_177 
* INOUT : bl_0_178 
* INOUT : br_0_178 
* INOUT : bl_0_179 
* INOUT : br_0_179 
* INOUT : bl_0_180 
* INOUT : br_0_180 
* INOUT : bl_0_181 
* INOUT : br_0_181 
* INOUT : bl_0_182 
* INOUT : br_0_182 
* INOUT : bl_0_183 
* INOUT : br_0_183 
* INOUT : bl_0_184 
* INOUT : br_0_184 
* INOUT : bl_0_185 
* INOUT : br_0_185 
* INOUT : bl_0_186 
* INOUT : br_0_186 
* INOUT : bl_0_187 
* INOUT : br_0_187 
* INOUT : bl_0_188 
* INOUT : br_0_188 
* INOUT : bl_0_189 
* INOUT : br_0_189 
* INOUT : bl_0_190 
* INOUT : br_0_190 
* INOUT : bl_0_191 
* INOUT : br_0_191 
* INOUT : bl_0_192 
* INOUT : br_0_192 
* INOUT : bl_0_193 
* INOUT : br_0_193 
* INOUT : bl_0_194 
* INOUT : br_0_194 
* INOUT : bl_0_195 
* INOUT : br_0_195 
* INOUT : bl_0_196 
* INOUT : br_0_196 
* INOUT : bl_0_197 
* INOUT : br_0_197 
* INOUT : bl_0_198 
* INOUT : br_0_198 
* INOUT : bl_0_199 
* INOUT : br_0_199 
* INOUT : bl_0_200 
* INOUT : br_0_200 
* INOUT : bl_0_201 
* INOUT : br_0_201 
* INOUT : bl_0_202 
* INOUT : br_0_202 
* INOUT : bl_0_203 
* INOUT : br_0_203 
* INOUT : bl_0_204 
* INOUT : br_0_204 
* INOUT : bl_0_205 
* INOUT : br_0_205 
* INOUT : bl_0_206 
* INOUT : br_0_206 
* INOUT : bl_0_207 
* INOUT : br_0_207 
* INOUT : bl_0_208 
* INOUT : br_0_208 
* INOUT : bl_0_209 
* INOUT : br_0_209 
* INOUT : bl_0_210 
* INOUT : br_0_210 
* INOUT : bl_0_211 
* INOUT : br_0_211 
* INOUT : bl_0_212 
* INOUT : br_0_212 
* INOUT : bl_0_213 
* INOUT : br_0_213 
* INOUT : bl_0_214 
* INOUT : br_0_214 
* INOUT : bl_0_215 
* INOUT : br_0_215 
* INOUT : bl_0_216 
* INOUT : br_0_216 
* INOUT : bl_0_217 
* INOUT : br_0_217 
* INOUT : bl_0_218 
* INOUT : br_0_218 
* INOUT : bl_0_219 
* INOUT : br_0_219 
* INOUT : bl_0_220 
* INOUT : br_0_220 
* INOUT : bl_0_221 
* INOUT : br_0_221 
* INOUT : bl_0_222 
* INOUT : br_0_222 
* INOUT : bl_0_223 
* INOUT : br_0_223 
* INOUT : bl_0_224 
* INOUT : br_0_224 
* INOUT : bl_0_225 
* INOUT : br_0_225 
* INOUT : bl_0_226 
* INOUT : br_0_226 
* INOUT : bl_0_227 
* INOUT : br_0_227 
* INOUT : bl_0_228 
* INOUT : br_0_228 
* INOUT : bl_0_229 
* INOUT : br_0_229 
* INOUT : bl_0_230 
* INOUT : br_0_230 
* INOUT : bl_0_231 
* INOUT : br_0_231 
* INOUT : bl_0_232 
* INOUT : br_0_232 
* INOUT : bl_0_233 
* INOUT : br_0_233 
* INOUT : bl_0_234 
* INOUT : br_0_234 
* INOUT : bl_0_235 
* INOUT : br_0_235 
* INOUT : bl_0_236 
* INOUT : br_0_236 
* INOUT : bl_0_237 
* INOUT : br_0_237 
* INOUT : bl_0_238 
* INOUT : br_0_238 
* INOUT : bl_0_239 
* INOUT : br_0_239 
* INOUT : bl_0_240 
* INOUT : br_0_240 
* INOUT : bl_0_241 
* INOUT : br_0_241 
* INOUT : bl_0_242 
* INOUT : br_0_242 
* INOUT : bl_0_243 
* INOUT : br_0_243 
* INOUT : bl_0_244 
* INOUT : br_0_244 
* INOUT : bl_0_245 
* INOUT : br_0_245 
* INOUT : bl_0_246 
* INOUT : br_0_246 
* INOUT : bl_0_247 
* INOUT : br_0_247 
* INOUT : bl_0_248 
* INOUT : br_0_248 
* INOUT : bl_0_249 
* INOUT : br_0_249 
* INOUT : bl_0_250 
* INOUT : br_0_250 
* INOUT : bl_0_251 
* INOUT : br_0_251 
* INOUT : bl_0_252 
* INOUT : br_0_252 
* INOUT : bl_0_253 
* INOUT : br_0_253 
* INOUT : bl_0_254 
* INOUT : br_0_254 
* INOUT : bl_0_255 
* INOUT : br_0_255 
* INPUT : rbl_wl_0_0 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* INPUT : wl_0_33 
* INPUT : wl_0_34 
* INPUT : wl_0_35 
* INPUT : wl_0_36 
* INPUT : wl_0_37 
* INPUT : wl_0_38 
* INPUT : wl_0_39 
* INPUT : wl_0_40 
* INPUT : wl_0_41 
* INPUT : wl_0_42 
* INPUT : wl_0_43 
* INPUT : wl_0_44 
* INPUT : wl_0_45 
* INPUT : wl_0_46 
* INPUT : wl_0_47 
* INPUT : wl_0_48 
* INPUT : wl_0_49 
* INPUT : wl_0_50 
* INPUT : wl_0_51 
* INPUT : wl_0_52 
* INPUT : wl_0_53 
* INPUT : wl_0_54 
* INPUT : wl_0_55 
* INPUT : wl_0_56 
* INPUT : wl_0_57 
* INPUT : wl_0_58 
* INPUT : wl_0_59 
* INPUT : wl_0_60 
* INPUT : wl_0_61 
* INPUT : wl_0_62 
* INPUT : wl_0_63 
* INPUT : wl_0_64 
* INPUT : wl_0_65 
* INPUT : wl_0_66 
* INPUT : wl_0_67 
* INPUT : wl_0_68 
* INPUT : wl_0_69 
* INPUT : wl_0_70 
* INPUT : wl_0_71 
* INPUT : wl_0_72 
* INPUT : wl_0_73 
* INPUT : wl_0_74 
* INPUT : wl_0_75 
* INPUT : wl_0_76 
* INPUT : wl_0_77 
* INPUT : wl_0_78 
* INPUT : wl_0_79 
* INPUT : wl_0_80 
* INPUT : wl_0_81 
* INPUT : wl_0_82 
* INPUT : wl_0_83 
* INPUT : wl_0_84 
* INPUT : wl_0_85 
* INPUT : wl_0_86 
* INPUT : wl_0_87 
* INPUT : wl_0_88 
* INPUT : wl_0_89 
* INPUT : wl_0_90 
* INPUT : wl_0_91 
* INPUT : wl_0_92 
* INPUT : wl_0_93 
* INPUT : wl_0_94 
* INPUT : wl_0_95 
* INPUT : wl_0_96 
* INPUT : wl_0_97 
* INPUT : wl_0_98 
* INPUT : wl_0_99 
* INPUT : wl_0_100 
* INPUT : wl_0_101 
* INPUT : wl_0_102 
* INPUT : wl_0_103 
* INPUT : wl_0_104 
* INPUT : wl_0_105 
* INPUT : wl_0_106 
* INPUT : wl_0_107 
* INPUT : wl_0_108 
* INPUT : wl_0_109 
* INPUT : wl_0_110 
* INPUT : wl_0_111 
* INPUT : wl_0_112 
* INPUT : wl_0_113 
* INPUT : wl_0_114 
* INPUT : wl_0_115 
* INPUT : wl_0_116 
* INPUT : wl_0_117 
* INPUT : wl_0_118 
* INPUT : wl_0_119 
* INPUT : wl_0_120 
* INPUT : wl_0_121 
* INPUT : wl_0_122 
* INPUT : wl_0_123 
* INPUT : wl_0_124 
* INPUT : wl_0_125 
* INPUT : wl_0_126 
* INPUT : wl_0_127 
* POWER : vdd 
* GROUND: gnd 
* rows: 128 cols: 256
* rbl: [1, 0] left_rbl: [0] right_rbl: []
Xbitcell_array
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65
+ bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69
+ bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73
+ bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77
+ bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81
+ bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85
+ bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89
+ bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93
+ bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97
+ bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101
+ bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105
+ br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108
+ bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112
+ br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115
+ bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119
+ br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122
+ bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126
+ br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 bl_0_129 br_0_129
+ bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132 br_0_132 bl_0_133
+ br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135 bl_0_136 br_0_136
+ bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139 br_0_139 bl_0_140
+ br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142 bl_0_143 br_0_143
+ bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146 br_0_146 bl_0_147
+ br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149 bl_0_150 br_0_150
+ bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153 br_0_153 bl_0_154
+ br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156 bl_0_157 br_0_157
+ bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160 br_0_160 bl_0_161
+ br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163 bl_0_164 br_0_164
+ bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167 br_0_167 bl_0_168
+ br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170 bl_0_171 br_0_171
+ bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174 br_0_174 bl_0_175
+ br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177 bl_0_178 br_0_178
+ bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181 br_0_181 bl_0_182
+ br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184 bl_0_185 br_0_185
+ bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188 br_0_188 bl_0_189
+ br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191 bl_0_192 br_0_192
+ bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195 br_0_195 bl_0_196
+ br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198 bl_0_199 br_0_199
+ bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202 br_0_202 bl_0_203
+ br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205 bl_0_206 br_0_206
+ bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209 br_0_209 bl_0_210
+ br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212 bl_0_213 br_0_213
+ bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216 br_0_216 bl_0_217
+ br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219 bl_0_220 br_0_220
+ bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223 br_0_223 bl_0_224
+ br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226 bl_0_227 br_0_227
+ bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230 br_0_230 bl_0_231
+ br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233 bl_0_234 br_0_234
+ bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237 br_0_237 bl_0_238
+ br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240 bl_0_241 br_0_241
+ bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244 br_0_244 bl_0_245
+ br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247 bl_0_248 br_0_248
+ bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251 br_0_251 bl_0_252
+ br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254 bl_0_255 br_0_255 wl_0_0
+ wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10
+ wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18
+ wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26
+ wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34
+ wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42
+ wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50
+ wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57 wl_0_58
+ wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 wl_0_65 wl_0_66
+ wl_0_67 wl_0_68 wl_0_69 wl_0_70 wl_0_71 wl_0_72 wl_0_73 wl_0_74
+ wl_0_75 wl_0_76 wl_0_77 wl_0_78 wl_0_79 wl_0_80 wl_0_81 wl_0_82
+ wl_0_83 wl_0_84 wl_0_85 wl_0_86 wl_0_87 wl_0_88 wl_0_89 wl_0_90
+ wl_0_91 wl_0_92 wl_0_93 wl_0_94 wl_0_95 wl_0_96 wl_0_97 wl_0_98
+ wl_0_99 wl_0_100 wl_0_101 wl_0_102 wl_0_103 wl_0_104 wl_0_105 wl_0_106
+ wl_0_107 wl_0_108 wl_0_109 wl_0_110 wl_0_111 wl_0_112 wl_0_113
+ wl_0_114 wl_0_115 wl_0_116 wl_0_117 wl_0_118 wl_0_119 wl_0_120
+ wl_0_121 wl_0_122 wl_0_123 wl_0_124 wl_0_125 wl_0_126 wl_0_127 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_bitcell_array
Xreplica_col_0
+ rbl_bl_0_0 rbl_br_0_0 rbl_wl_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4
+ wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13
+ wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21
+ wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29
+ wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37
+ wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45
+ wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53
+ wl_0_54 wl_0_55 wl_0_56 wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61
+ wl_0_62 wl_0_63 wl_0_64 wl_0_65 wl_0_66 wl_0_67 wl_0_68 wl_0_69
+ wl_0_70 wl_0_71 wl_0_72 wl_0_73 wl_0_74 wl_0_75 wl_0_76 wl_0_77
+ wl_0_78 wl_0_79 wl_0_80 wl_0_81 wl_0_82 wl_0_83 wl_0_84 wl_0_85
+ wl_0_86 wl_0_87 wl_0_88 wl_0_89 wl_0_90 wl_0_91 wl_0_92 wl_0_93
+ wl_0_94 wl_0_95 wl_0_96 wl_0_97 wl_0_98 wl_0_99 wl_0_100 wl_0_101
+ wl_0_102 wl_0_103 wl_0_104 wl_0_105 wl_0_106 wl_0_107 wl_0_108
+ wl_0_109 wl_0_110 wl_0_111 wl_0_112 wl_0_113 wl_0_114 wl_0_115
+ wl_0_116 wl_0_117 wl_0_118 wl_0_119 wl_0_120 wl_0_121 wl_0_122
+ wl_0_123 wl_0_124 wl_0_125 wl_0_126 wl_0_127 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_replica_column
Xdummy_row_0
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65
+ bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69
+ bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73
+ bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77
+ bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81
+ bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85
+ bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89
+ bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93
+ bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97
+ bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101
+ bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105
+ br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108
+ bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112
+ br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115
+ bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119
+ br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122
+ bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126
+ br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 bl_0_129 br_0_129
+ bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132 br_0_132 bl_0_133
+ br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135 bl_0_136 br_0_136
+ bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139 br_0_139 bl_0_140
+ br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142 bl_0_143 br_0_143
+ bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146 br_0_146 bl_0_147
+ br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149 bl_0_150 br_0_150
+ bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153 br_0_153 bl_0_154
+ br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156 bl_0_157 br_0_157
+ bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160 br_0_160 bl_0_161
+ br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163 bl_0_164 br_0_164
+ bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167 br_0_167 bl_0_168
+ br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170 bl_0_171 br_0_171
+ bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174 br_0_174 bl_0_175
+ br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177 bl_0_178 br_0_178
+ bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181 br_0_181 bl_0_182
+ br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184 bl_0_185 br_0_185
+ bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188 br_0_188 bl_0_189
+ br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191 bl_0_192 br_0_192
+ bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195 br_0_195 bl_0_196
+ br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198 bl_0_199 br_0_199
+ bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202 br_0_202 bl_0_203
+ br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205 bl_0_206 br_0_206
+ bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209 br_0_209 bl_0_210
+ br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212 bl_0_213 br_0_213
+ bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216 br_0_216 bl_0_217
+ br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219 bl_0_220 br_0_220
+ bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223 br_0_223 bl_0_224
+ br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226 bl_0_227 br_0_227
+ bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230 br_0_230 bl_0_231
+ br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233 bl_0_234 br_0_234
+ bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237 br_0_237 bl_0_238
+ br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240 bl_0_241 br_0_241
+ bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244 br_0_244 bl_0_245
+ br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247 bl_0_248 br_0_248
+ bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251 br_0_251 bl_0_252
+ br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254 bl_0_255 br_0_255
+ rbl_wl_0_0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_dummy_array
.ENDS sram_1rw0r0w_32_1024_freepdk45_replica_bitcell_array

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_dummy_array_2
+ bl_0_0 br_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7
+ wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16
+ wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24
+ wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32
+ wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40
+ wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48
+ wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56
+ wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64
+ wl_0_65 wl_0_66 wl_0_67 wl_0_68 wl_0_69 wl_0_70 wl_0_71 wl_0_72
+ wl_0_73 wl_0_74 wl_0_75 wl_0_76 wl_0_77 wl_0_78 wl_0_79 wl_0_80
+ wl_0_81 wl_0_82 wl_0_83 wl_0_84 wl_0_85 wl_0_86 wl_0_87 wl_0_88
+ wl_0_89 wl_0_90 wl_0_91 wl_0_92 wl_0_93 wl_0_94 wl_0_95 wl_0_96
+ wl_0_97 wl_0_98 wl_0_99 wl_0_100 wl_0_101 wl_0_102 wl_0_103 wl_0_104
+ wl_0_105 wl_0_106 wl_0_107 wl_0_108 wl_0_109 wl_0_110 wl_0_111
+ wl_0_112 wl_0_113 wl_0_114 wl_0_115 wl_0_116 wl_0_117 wl_0_118
+ wl_0_119 wl_0_120 wl_0_121 wl_0_122 wl_0_123 wl_0_124 wl_0_125
+ wl_0_126 wl_0_127 wl_0_128 wl_0_129 wl_0_130 vdd gnd
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* INPUT : wl_0_33 
* INPUT : wl_0_34 
* INPUT : wl_0_35 
* INPUT : wl_0_36 
* INPUT : wl_0_37 
* INPUT : wl_0_38 
* INPUT : wl_0_39 
* INPUT : wl_0_40 
* INPUT : wl_0_41 
* INPUT : wl_0_42 
* INPUT : wl_0_43 
* INPUT : wl_0_44 
* INPUT : wl_0_45 
* INPUT : wl_0_46 
* INPUT : wl_0_47 
* INPUT : wl_0_48 
* INPUT : wl_0_49 
* INPUT : wl_0_50 
* INPUT : wl_0_51 
* INPUT : wl_0_52 
* INPUT : wl_0_53 
* INPUT : wl_0_54 
* INPUT : wl_0_55 
* INPUT : wl_0_56 
* INPUT : wl_0_57 
* INPUT : wl_0_58 
* INPUT : wl_0_59 
* INPUT : wl_0_60 
* INPUT : wl_0_61 
* INPUT : wl_0_62 
* INPUT : wl_0_63 
* INPUT : wl_0_64 
* INPUT : wl_0_65 
* INPUT : wl_0_66 
* INPUT : wl_0_67 
* INPUT : wl_0_68 
* INPUT : wl_0_69 
* INPUT : wl_0_70 
* INPUT : wl_0_71 
* INPUT : wl_0_72 
* INPUT : wl_0_73 
* INPUT : wl_0_74 
* INPUT : wl_0_75 
* INPUT : wl_0_76 
* INPUT : wl_0_77 
* INPUT : wl_0_78 
* INPUT : wl_0_79 
* INPUT : wl_0_80 
* INPUT : wl_0_81 
* INPUT : wl_0_82 
* INPUT : wl_0_83 
* INPUT : wl_0_84 
* INPUT : wl_0_85 
* INPUT : wl_0_86 
* INPUT : wl_0_87 
* INPUT : wl_0_88 
* INPUT : wl_0_89 
* INPUT : wl_0_90 
* INPUT : wl_0_91 
* INPUT : wl_0_92 
* INPUT : wl_0_93 
* INPUT : wl_0_94 
* INPUT : wl_0_95 
* INPUT : wl_0_96 
* INPUT : wl_0_97 
* INPUT : wl_0_98 
* INPUT : wl_0_99 
* INPUT : wl_0_100 
* INPUT : wl_0_101 
* INPUT : wl_0_102 
* INPUT : wl_0_103 
* INPUT : wl_0_104 
* INPUT : wl_0_105 
* INPUT : wl_0_106 
* INPUT : wl_0_107 
* INPUT : wl_0_108 
* INPUT : wl_0_109 
* INPUT : wl_0_110 
* INPUT : wl_0_111 
* INPUT : wl_0_112 
* INPUT : wl_0_113 
* INPUT : wl_0_114 
* INPUT : wl_0_115 
* INPUT : wl_0_116 
* INPUT : wl_0_117 
* INPUT : wl_0_118 
* INPUT : wl_0_119 
* INPUT : wl_0_120 
* INPUT : wl_0_121 
* INPUT : wl_0_122 
* INPUT : wl_0_123 
* INPUT : wl_0_124 
* INPUT : wl_0_125 
* INPUT : wl_0_126 
* INPUT : wl_0_127 
* INPUT : wl_0_128 
* INPUT : wl_0_129 
* INPUT : wl_0_130 
* POWER : vdd 
* GROUND: gnd 
Xbit_r0_c0
+ bl_0_0 br_0_0 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r1_c0
+ bl_0_0 br_0_0 wl_0_1 vdd gnd
+ dummy_cell_1rw
Xbit_r2_c0
+ bl_0_0 br_0_0 wl_0_2 vdd gnd
+ dummy_cell_1rw
Xbit_r3_c0
+ bl_0_0 br_0_0 wl_0_3 vdd gnd
+ dummy_cell_1rw
Xbit_r4_c0
+ bl_0_0 br_0_0 wl_0_4 vdd gnd
+ dummy_cell_1rw
Xbit_r5_c0
+ bl_0_0 br_0_0 wl_0_5 vdd gnd
+ dummy_cell_1rw
Xbit_r6_c0
+ bl_0_0 br_0_0 wl_0_6 vdd gnd
+ dummy_cell_1rw
Xbit_r7_c0
+ bl_0_0 br_0_0 wl_0_7 vdd gnd
+ dummy_cell_1rw
Xbit_r8_c0
+ bl_0_0 br_0_0 wl_0_8 vdd gnd
+ dummy_cell_1rw
Xbit_r9_c0
+ bl_0_0 br_0_0 wl_0_9 vdd gnd
+ dummy_cell_1rw
Xbit_r10_c0
+ bl_0_0 br_0_0 wl_0_10 vdd gnd
+ dummy_cell_1rw
Xbit_r11_c0
+ bl_0_0 br_0_0 wl_0_11 vdd gnd
+ dummy_cell_1rw
Xbit_r12_c0
+ bl_0_0 br_0_0 wl_0_12 vdd gnd
+ dummy_cell_1rw
Xbit_r13_c0
+ bl_0_0 br_0_0 wl_0_13 vdd gnd
+ dummy_cell_1rw
Xbit_r14_c0
+ bl_0_0 br_0_0 wl_0_14 vdd gnd
+ dummy_cell_1rw
Xbit_r15_c0
+ bl_0_0 br_0_0 wl_0_15 vdd gnd
+ dummy_cell_1rw
Xbit_r16_c0
+ bl_0_0 br_0_0 wl_0_16 vdd gnd
+ dummy_cell_1rw
Xbit_r17_c0
+ bl_0_0 br_0_0 wl_0_17 vdd gnd
+ dummy_cell_1rw
Xbit_r18_c0
+ bl_0_0 br_0_0 wl_0_18 vdd gnd
+ dummy_cell_1rw
Xbit_r19_c0
+ bl_0_0 br_0_0 wl_0_19 vdd gnd
+ dummy_cell_1rw
Xbit_r20_c0
+ bl_0_0 br_0_0 wl_0_20 vdd gnd
+ dummy_cell_1rw
Xbit_r21_c0
+ bl_0_0 br_0_0 wl_0_21 vdd gnd
+ dummy_cell_1rw
Xbit_r22_c0
+ bl_0_0 br_0_0 wl_0_22 vdd gnd
+ dummy_cell_1rw
Xbit_r23_c0
+ bl_0_0 br_0_0 wl_0_23 vdd gnd
+ dummy_cell_1rw
Xbit_r24_c0
+ bl_0_0 br_0_0 wl_0_24 vdd gnd
+ dummy_cell_1rw
Xbit_r25_c0
+ bl_0_0 br_0_0 wl_0_25 vdd gnd
+ dummy_cell_1rw
Xbit_r26_c0
+ bl_0_0 br_0_0 wl_0_26 vdd gnd
+ dummy_cell_1rw
Xbit_r27_c0
+ bl_0_0 br_0_0 wl_0_27 vdd gnd
+ dummy_cell_1rw
Xbit_r28_c0
+ bl_0_0 br_0_0 wl_0_28 vdd gnd
+ dummy_cell_1rw
Xbit_r29_c0
+ bl_0_0 br_0_0 wl_0_29 vdd gnd
+ dummy_cell_1rw
Xbit_r30_c0
+ bl_0_0 br_0_0 wl_0_30 vdd gnd
+ dummy_cell_1rw
Xbit_r31_c0
+ bl_0_0 br_0_0 wl_0_31 vdd gnd
+ dummy_cell_1rw
Xbit_r32_c0
+ bl_0_0 br_0_0 wl_0_32 vdd gnd
+ dummy_cell_1rw
Xbit_r33_c0
+ bl_0_0 br_0_0 wl_0_33 vdd gnd
+ dummy_cell_1rw
Xbit_r34_c0
+ bl_0_0 br_0_0 wl_0_34 vdd gnd
+ dummy_cell_1rw
Xbit_r35_c0
+ bl_0_0 br_0_0 wl_0_35 vdd gnd
+ dummy_cell_1rw
Xbit_r36_c0
+ bl_0_0 br_0_0 wl_0_36 vdd gnd
+ dummy_cell_1rw
Xbit_r37_c0
+ bl_0_0 br_0_0 wl_0_37 vdd gnd
+ dummy_cell_1rw
Xbit_r38_c0
+ bl_0_0 br_0_0 wl_0_38 vdd gnd
+ dummy_cell_1rw
Xbit_r39_c0
+ bl_0_0 br_0_0 wl_0_39 vdd gnd
+ dummy_cell_1rw
Xbit_r40_c0
+ bl_0_0 br_0_0 wl_0_40 vdd gnd
+ dummy_cell_1rw
Xbit_r41_c0
+ bl_0_0 br_0_0 wl_0_41 vdd gnd
+ dummy_cell_1rw
Xbit_r42_c0
+ bl_0_0 br_0_0 wl_0_42 vdd gnd
+ dummy_cell_1rw
Xbit_r43_c0
+ bl_0_0 br_0_0 wl_0_43 vdd gnd
+ dummy_cell_1rw
Xbit_r44_c0
+ bl_0_0 br_0_0 wl_0_44 vdd gnd
+ dummy_cell_1rw
Xbit_r45_c0
+ bl_0_0 br_0_0 wl_0_45 vdd gnd
+ dummy_cell_1rw
Xbit_r46_c0
+ bl_0_0 br_0_0 wl_0_46 vdd gnd
+ dummy_cell_1rw
Xbit_r47_c0
+ bl_0_0 br_0_0 wl_0_47 vdd gnd
+ dummy_cell_1rw
Xbit_r48_c0
+ bl_0_0 br_0_0 wl_0_48 vdd gnd
+ dummy_cell_1rw
Xbit_r49_c0
+ bl_0_0 br_0_0 wl_0_49 vdd gnd
+ dummy_cell_1rw
Xbit_r50_c0
+ bl_0_0 br_0_0 wl_0_50 vdd gnd
+ dummy_cell_1rw
Xbit_r51_c0
+ bl_0_0 br_0_0 wl_0_51 vdd gnd
+ dummy_cell_1rw
Xbit_r52_c0
+ bl_0_0 br_0_0 wl_0_52 vdd gnd
+ dummy_cell_1rw
Xbit_r53_c0
+ bl_0_0 br_0_0 wl_0_53 vdd gnd
+ dummy_cell_1rw
Xbit_r54_c0
+ bl_0_0 br_0_0 wl_0_54 vdd gnd
+ dummy_cell_1rw
Xbit_r55_c0
+ bl_0_0 br_0_0 wl_0_55 vdd gnd
+ dummy_cell_1rw
Xbit_r56_c0
+ bl_0_0 br_0_0 wl_0_56 vdd gnd
+ dummy_cell_1rw
Xbit_r57_c0
+ bl_0_0 br_0_0 wl_0_57 vdd gnd
+ dummy_cell_1rw
Xbit_r58_c0
+ bl_0_0 br_0_0 wl_0_58 vdd gnd
+ dummy_cell_1rw
Xbit_r59_c0
+ bl_0_0 br_0_0 wl_0_59 vdd gnd
+ dummy_cell_1rw
Xbit_r60_c0
+ bl_0_0 br_0_0 wl_0_60 vdd gnd
+ dummy_cell_1rw
Xbit_r61_c0
+ bl_0_0 br_0_0 wl_0_61 vdd gnd
+ dummy_cell_1rw
Xbit_r62_c0
+ bl_0_0 br_0_0 wl_0_62 vdd gnd
+ dummy_cell_1rw
Xbit_r63_c0
+ bl_0_0 br_0_0 wl_0_63 vdd gnd
+ dummy_cell_1rw
Xbit_r64_c0
+ bl_0_0 br_0_0 wl_0_64 vdd gnd
+ dummy_cell_1rw
Xbit_r65_c0
+ bl_0_0 br_0_0 wl_0_65 vdd gnd
+ dummy_cell_1rw
Xbit_r66_c0
+ bl_0_0 br_0_0 wl_0_66 vdd gnd
+ dummy_cell_1rw
Xbit_r67_c0
+ bl_0_0 br_0_0 wl_0_67 vdd gnd
+ dummy_cell_1rw
Xbit_r68_c0
+ bl_0_0 br_0_0 wl_0_68 vdd gnd
+ dummy_cell_1rw
Xbit_r69_c0
+ bl_0_0 br_0_0 wl_0_69 vdd gnd
+ dummy_cell_1rw
Xbit_r70_c0
+ bl_0_0 br_0_0 wl_0_70 vdd gnd
+ dummy_cell_1rw
Xbit_r71_c0
+ bl_0_0 br_0_0 wl_0_71 vdd gnd
+ dummy_cell_1rw
Xbit_r72_c0
+ bl_0_0 br_0_0 wl_0_72 vdd gnd
+ dummy_cell_1rw
Xbit_r73_c0
+ bl_0_0 br_0_0 wl_0_73 vdd gnd
+ dummy_cell_1rw
Xbit_r74_c0
+ bl_0_0 br_0_0 wl_0_74 vdd gnd
+ dummy_cell_1rw
Xbit_r75_c0
+ bl_0_0 br_0_0 wl_0_75 vdd gnd
+ dummy_cell_1rw
Xbit_r76_c0
+ bl_0_0 br_0_0 wl_0_76 vdd gnd
+ dummy_cell_1rw
Xbit_r77_c0
+ bl_0_0 br_0_0 wl_0_77 vdd gnd
+ dummy_cell_1rw
Xbit_r78_c0
+ bl_0_0 br_0_0 wl_0_78 vdd gnd
+ dummy_cell_1rw
Xbit_r79_c0
+ bl_0_0 br_0_0 wl_0_79 vdd gnd
+ dummy_cell_1rw
Xbit_r80_c0
+ bl_0_0 br_0_0 wl_0_80 vdd gnd
+ dummy_cell_1rw
Xbit_r81_c0
+ bl_0_0 br_0_0 wl_0_81 vdd gnd
+ dummy_cell_1rw
Xbit_r82_c0
+ bl_0_0 br_0_0 wl_0_82 vdd gnd
+ dummy_cell_1rw
Xbit_r83_c0
+ bl_0_0 br_0_0 wl_0_83 vdd gnd
+ dummy_cell_1rw
Xbit_r84_c0
+ bl_0_0 br_0_0 wl_0_84 vdd gnd
+ dummy_cell_1rw
Xbit_r85_c0
+ bl_0_0 br_0_0 wl_0_85 vdd gnd
+ dummy_cell_1rw
Xbit_r86_c0
+ bl_0_0 br_0_0 wl_0_86 vdd gnd
+ dummy_cell_1rw
Xbit_r87_c0
+ bl_0_0 br_0_0 wl_0_87 vdd gnd
+ dummy_cell_1rw
Xbit_r88_c0
+ bl_0_0 br_0_0 wl_0_88 vdd gnd
+ dummy_cell_1rw
Xbit_r89_c0
+ bl_0_0 br_0_0 wl_0_89 vdd gnd
+ dummy_cell_1rw
Xbit_r90_c0
+ bl_0_0 br_0_0 wl_0_90 vdd gnd
+ dummy_cell_1rw
Xbit_r91_c0
+ bl_0_0 br_0_0 wl_0_91 vdd gnd
+ dummy_cell_1rw
Xbit_r92_c0
+ bl_0_0 br_0_0 wl_0_92 vdd gnd
+ dummy_cell_1rw
Xbit_r93_c0
+ bl_0_0 br_0_0 wl_0_93 vdd gnd
+ dummy_cell_1rw
Xbit_r94_c0
+ bl_0_0 br_0_0 wl_0_94 vdd gnd
+ dummy_cell_1rw
Xbit_r95_c0
+ bl_0_0 br_0_0 wl_0_95 vdd gnd
+ dummy_cell_1rw
Xbit_r96_c0
+ bl_0_0 br_0_0 wl_0_96 vdd gnd
+ dummy_cell_1rw
Xbit_r97_c0
+ bl_0_0 br_0_0 wl_0_97 vdd gnd
+ dummy_cell_1rw
Xbit_r98_c0
+ bl_0_0 br_0_0 wl_0_98 vdd gnd
+ dummy_cell_1rw
Xbit_r99_c0
+ bl_0_0 br_0_0 wl_0_99 vdd gnd
+ dummy_cell_1rw
Xbit_r100_c0
+ bl_0_0 br_0_0 wl_0_100 vdd gnd
+ dummy_cell_1rw
Xbit_r101_c0
+ bl_0_0 br_0_0 wl_0_101 vdd gnd
+ dummy_cell_1rw
Xbit_r102_c0
+ bl_0_0 br_0_0 wl_0_102 vdd gnd
+ dummy_cell_1rw
Xbit_r103_c0
+ bl_0_0 br_0_0 wl_0_103 vdd gnd
+ dummy_cell_1rw
Xbit_r104_c0
+ bl_0_0 br_0_0 wl_0_104 vdd gnd
+ dummy_cell_1rw
Xbit_r105_c0
+ bl_0_0 br_0_0 wl_0_105 vdd gnd
+ dummy_cell_1rw
Xbit_r106_c0
+ bl_0_0 br_0_0 wl_0_106 vdd gnd
+ dummy_cell_1rw
Xbit_r107_c0
+ bl_0_0 br_0_0 wl_0_107 vdd gnd
+ dummy_cell_1rw
Xbit_r108_c0
+ bl_0_0 br_0_0 wl_0_108 vdd gnd
+ dummy_cell_1rw
Xbit_r109_c0
+ bl_0_0 br_0_0 wl_0_109 vdd gnd
+ dummy_cell_1rw
Xbit_r110_c0
+ bl_0_0 br_0_0 wl_0_110 vdd gnd
+ dummy_cell_1rw
Xbit_r111_c0
+ bl_0_0 br_0_0 wl_0_111 vdd gnd
+ dummy_cell_1rw
Xbit_r112_c0
+ bl_0_0 br_0_0 wl_0_112 vdd gnd
+ dummy_cell_1rw
Xbit_r113_c0
+ bl_0_0 br_0_0 wl_0_113 vdd gnd
+ dummy_cell_1rw
Xbit_r114_c0
+ bl_0_0 br_0_0 wl_0_114 vdd gnd
+ dummy_cell_1rw
Xbit_r115_c0
+ bl_0_0 br_0_0 wl_0_115 vdd gnd
+ dummy_cell_1rw
Xbit_r116_c0
+ bl_0_0 br_0_0 wl_0_116 vdd gnd
+ dummy_cell_1rw
Xbit_r117_c0
+ bl_0_0 br_0_0 wl_0_117 vdd gnd
+ dummy_cell_1rw
Xbit_r118_c0
+ bl_0_0 br_0_0 wl_0_118 vdd gnd
+ dummy_cell_1rw
Xbit_r119_c0
+ bl_0_0 br_0_0 wl_0_119 vdd gnd
+ dummy_cell_1rw
Xbit_r120_c0
+ bl_0_0 br_0_0 wl_0_120 vdd gnd
+ dummy_cell_1rw
Xbit_r121_c0
+ bl_0_0 br_0_0 wl_0_121 vdd gnd
+ dummy_cell_1rw
Xbit_r122_c0
+ bl_0_0 br_0_0 wl_0_122 vdd gnd
+ dummy_cell_1rw
Xbit_r123_c0
+ bl_0_0 br_0_0 wl_0_123 vdd gnd
+ dummy_cell_1rw
Xbit_r124_c0
+ bl_0_0 br_0_0 wl_0_124 vdd gnd
+ dummy_cell_1rw
Xbit_r125_c0
+ bl_0_0 br_0_0 wl_0_125 vdd gnd
+ dummy_cell_1rw
Xbit_r126_c0
+ bl_0_0 br_0_0 wl_0_126 vdd gnd
+ dummy_cell_1rw
Xbit_r127_c0
+ bl_0_0 br_0_0 wl_0_127 vdd gnd
+ dummy_cell_1rw
Xbit_r128_c0
+ bl_0_0 br_0_0 wl_0_128 vdd gnd
+ dummy_cell_1rw
Xbit_r129_c0
+ bl_0_0 br_0_0 wl_0_129 vdd gnd
+ dummy_cell_1rw
Xbit_r130_c0
+ bl_0_0 br_0_0 wl_0_130 vdd gnd
+ dummy_cell_1rw
.ENDS sram_1rw0r0w_32_1024_freepdk45_dummy_array_2

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_dummy_array_0
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65
+ bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69
+ bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73
+ bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77
+ bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81
+ bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85
+ bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89
+ bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93
+ bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97
+ bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101
+ bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105
+ br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108
+ bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112
+ br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115
+ bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119
+ br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122
+ bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126
+ br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 bl_0_129 br_0_129
+ bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132 br_0_132 bl_0_133
+ br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135 bl_0_136 br_0_136
+ bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139 br_0_139 bl_0_140
+ br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142 bl_0_143 br_0_143
+ bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146 br_0_146 bl_0_147
+ br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149 bl_0_150 br_0_150
+ bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153 br_0_153 bl_0_154
+ br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156 bl_0_157 br_0_157
+ bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160 br_0_160 bl_0_161
+ br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163 bl_0_164 br_0_164
+ bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167 br_0_167 bl_0_168
+ br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170 bl_0_171 br_0_171
+ bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174 br_0_174 bl_0_175
+ br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177 bl_0_178 br_0_178
+ bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181 br_0_181 bl_0_182
+ br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184 bl_0_185 br_0_185
+ bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188 br_0_188 bl_0_189
+ br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191 bl_0_192 br_0_192
+ bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195 br_0_195 bl_0_196
+ br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198 bl_0_199 br_0_199
+ bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202 br_0_202 bl_0_203
+ br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205 bl_0_206 br_0_206
+ bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209 br_0_209 bl_0_210
+ br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212 bl_0_213 br_0_213
+ bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216 br_0_216 bl_0_217
+ br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219 bl_0_220 br_0_220
+ bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223 br_0_223 bl_0_224
+ br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226 bl_0_227 br_0_227
+ bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230 br_0_230 bl_0_231
+ br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233 bl_0_234 br_0_234
+ bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237 br_0_237 bl_0_238
+ br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240 bl_0_241 br_0_241
+ bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244 br_0_244 bl_0_245
+ br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247 bl_0_248 br_0_248
+ bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251 br_0_251 bl_0_252
+ br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254 bl_0_255 br_0_255
+ bl_0_256 br_0_256 wl_0_0 vdd gnd
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INOUT : bl_0_64 
* INOUT : br_0_64 
* INOUT : bl_0_65 
* INOUT : br_0_65 
* INOUT : bl_0_66 
* INOUT : br_0_66 
* INOUT : bl_0_67 
* INOUT : br_0_67 
* INOUT : bl_0_68 
* INOUT : br_0_68 
* INOUT : bl_0_69 
* INOUT : br_0_69 
* INOUT : bl_0_70 
* INOUT : br_0_70 
* INOUT : bl_0_71 
* INOUT : br_0_71 
* INOUT : bl_0_72 
* INOUT : br_0_72 
* INOUT : bl_0_73 
* INOUT : br_0_73 
* INOUT : bl_0_74 
* INOUT : br_0_74 
* INOUT : bl_0_75 
* INOUT : br_0_75 
* INOUT : bl_0_76 
* INOUT : br_0_76 
* INOUT : bl_0_77 
* INOUT : br_0_77 
* INOUT : bl_0_78 
* INOUT : br_0_78 
* INOUT : bl_0_79 
* INOUT : br_0_79 
* INOUT : bl_0_80 
* INOUT : br_0_80 
* INOUT : bl_0_81 
* INOUT : br_0_81 
* INOUT : bl_0_82 
* INOUT : br_0_82 
* INOUT : bl_0_83 
* INOUT : br_0_83 
* INOUT : bl_0_84 
* INOUT : br_0_84 
* INOUT : bl_0_85 
* INOUT : br_0_85 
* INOUT : bl_0_86 
* INOUT : br_0_86 
* INOUT : bl_0_87 
* INOUT : br_0_87 
* INOUT : bl_0_88 
* INOUT : br_0_88 
* INOUT : bl_0_89 
* INOUT : br_0_89 
* INOUT : bl_0_90 
* INOUT : br_0_90 
* INOUT : bl_0_91 
* INOUT : br_0_91 
* INOUT : bl_0_92 
* INOUT : br_0_92 
* INOUT : bl_0_93 
* INOUT : br_0_93 
* INOUT : bl_0_94 
* INOUT : br_0_94 
* INOUT : bl_0_95 
* INOUT : br_0_95 
* INOUT : bl_0_96 
* INOUT : br_0_96 
* INOUT : bl_0_97 
* INOUT : br_0_97 
* INOUT : bl_0_98 
* INOUT : br_0_98 
* INOUT : bl_0_99 
* INOUT : br_0_99 
* INOUT : bl_0_100 
* INOUT : br_0_100 
* INOUT : bl_0_101 
* INOUT : br_0_101 
* INOUT : bl_0_102 
* INOUT : br_0_102 
* INOUT : bl_0_103 
* INOUT : br_0_103 
* INOUT : bl_0_104 
* INOUT : br_0_104 
* INOUT : bl_0_105 
* INOUT : br_0_105 
* INOUT : bl_0_106 
* INOUT : br_0_106 
* INOUT : bl_0_107 
* INOUT : br_0_107 
* INOUT : bl_0_108 
* INOUT : br_0_108 
* INOUT : bl_0_109 
* INOUT : br_0_109 
* INOUT : bl_0_110 
* INOUT : br_0_110 
* INOUT : bl_0_111 
* INOUT : br_0_111 
* INOUT : bl_0_112 
* INOUT : br_0_112 
* INOUT : bl_0_113 
* INOUT : br_0_113 
* INOUT : bl_0_114 
* INOUT : br_0_114 
* INOUT : bl_0_115 
* INOUT : br_0_115 
* INOUT : bl_0_116 
* INOUT : br_0_116 
* INOUT : bl_0_117 
* INOUT : br_0_117 
* INOUT : bl_0_118 
* INOUT : br_0_118 
* INOUT : bl_0_119 
* INOUT : br_0_119 
* INOUT : bl_0_120 
* INOUT : br_0_120 
* INOUT : bl_0_121 
* INOUT : br_0_121 
* INOUT : bl_0_122 
* INOUT : br_0_122 
* INOUT : bl_0_123 
* INOUT : br_0_123 
* INOUT : bl_0_124 
* INOUT : br_0_124 
* INOUT : bl_0_125 
* INOUT : br_0_125 
* INOUT : bl_0_126 
* INOUT : br_0_126 
* INOUT : bl_0_127 
* INOUT : br_0_127 
* INOUT : bl_0_128 
* INOUT : br_0_128 
* INOUT : bl_0_129 
* INOUT : br_0_129 
* INOUT : bl_0_130 
* INOUT : br_0_130 
* INOUT : bl_0_131 
* INOUT : br_0_131 
* INOUT : bl_0_132 
* INOUT : br_0_132 
* INOUT : bl_0_133 
* INOUT : br_0_133 
* INOUT : bl_0_134 
* INOUT : br_0_134 
* INOUT : bl_0_135 
* INOUT : br_0_135 
* INOUT : bl_0_136 
* INOUT : br_0_136 
* INOUT : bl_0_137 
* INOUT : br_0_137 
* INOUT : bl_0_138 
* INOUT : br_0_138 
* INOUT : bl_0_139 
* INOUT : br_0_139 
* INOUT : bl_0_140 
* INOUT : br_0_140 
* INOUT : bl_0_141 
* INOUT : br_0_141 
* INOUT : bl_0_142 
* INOUT : br_0_142 
* INOUT : bl_0_143 
* INOUT : br_0_143 
* INOUT : bl_0_144 
* INOUT : br_0_144 
* INOUT : bl_0_145 
* INOUT : br_0_145 
* INOUT : bl_0_146 
* INOUT : br_0_146 
* INOUT : bl_0_147 
* INOUT : br_0_147 
* INOUT : bl_0_148 
* INOUT : br_0_148 
* INOUT : bl_0_149 
* INOUT : br_0_149 
* INOUT : bl_0_150 
* INOUT : br_0_150 
* INOUT : bl_0_151 
* INOUT : br_0_151 
* INOUT : bl_0_152 
* INOUT : br_0_152 
* INOUT : bl_0_153 
* INOUT : br_0_153 
* INOUT : bl_0_154 
* INOUT : br_0_154 
* INOUT : bl_0_155 
* INOUT : br_0_155 
* INOUT : bl_0_156 
* INOUT : br_0_156 
* INOUT : bl_0_157 
* INOUT : br_0_157 
* INOUT : bl_0_158 
* INOUT : br_0_158 
* INOUT : bl_0_159 
* INOUT : br_0_159 
* INOUT : bl_0_160 
* INOUT : br_0_160 
* INOUT : bl_0_161 
* INOUT : br_0_161 
* INOUT : bl_0_162 
* INOUT : br_0_162 
* INOUT : bl_0_163 
* INOUT : br_0_163 
* INOUT : bl_0_164 
* INOUT : br_0_164 
* INOUT : bl_0_165 
* INOUT : br_0_165 
* INOUT : bl_0_166 
* INOUT : br_0_166 
* INOUT : bl_0_167 
* INOUT : br_0_167 
* INOUT : bl_0_168 
* INOUT : br_0_168 
* INOUT : bl_0_169 
* INOUT : br_0_169 
* INOUT : bl_0_170 
* INOUT : br_0_170 
* INOUT : bl_0_171 
* INOUT : br_0_171 
* INOUT : bl_0_172 
* INOUT : br_0_172 
* INOUT : bl_0_173 
* INOUT : br_0_173 
* INOUT : bl_0_174 
* INOUT : br_0_174 
* INOUT : bl_0_175 
* INOUT : br_0_175 
* INOUT : bl_0_176 
* INOUT : br_0_176 
* INOUT : bl_0_177 
* INOUT : br_0_177 
* INOUT : bl_0_178 
* INOUT : br_0_178 
* INOUT : bl_0_179 
* INOUT : br_0_179 
* INOUT : bl_0_180 
* INOUT : br_0_180 
* INOUT : bl_0_181 
* INOUT : br_0_181 
* INOUT : bl_0_182 
* INOUT : br_0_182 
* INOUT : bl_0_183 
* INOUT : br_0_183 
* INOUT : bl_0_184 
* INOUT : br_0_184 
* INOUT : bl_0_185 
* INOUT : br_0_185 
* INOUT : bl_0_186 
* INOUT : br_0_186 
* INOUT : bl_0_187 
* INOUT : br_0_187 
* INOUT : bl_0_188 
* INOUT : br_0_188 
* INOUT : bl_0_189 
* INOUT : br_0_189 
* INOUT : bl_0_190 
* INOUT : br_0_190 
* INOUT : bl_0_191 
* INOUT : br_0_191 
* INOUT : bl_0_192 
* INOUT : br_0_192 
* INOUT : bl_0_193 
* INOUT : br_0_193 
* INOUT : bl_0_194 
* INOUT : br_0_194 
* INOUT : bl_0_195 
* INOUT : br_0_195 
* INOUT : bl_0_196 
* INOUT : br_0_196 
* INOUT : bl_0_197 
* INOUT : br_0_197 
* INOUT : bl_0_198 
* INOUT : br_0_198 
* INOUT : bl_0_199 
* INOUT : br_0_199 
* INOUT : bl_0_200 
* INOUT : br_0_200 
* INOUT : bl_0_201 
* INOUT : br_0_201 
* INOUT : bl_0_202 
* INOUT : br_0_202 
* INOUT : bl_0_203 
* INOUT : br_0_203 
* INOUT : bl_0_204 
* INOUT : br_0_204 
* INOUT : bl_0_205 
* INOUT : br_0_205 
* INOUT : bl_0_206 
* INOUT : br_0_206 
* INOUT : bl_0_207 
* INOUT : br_0_207 
* INOUT : bl_0_208 
* INOUT : br_0_208 
* INOUT : bl_0_209 
* INOUT : br_0_209 
* INOUT : bl_0_210 
* INOUT : br_0_210 
* INOUT : bl_0_211 
* INOUT : br_0_211 
* INOUT : bl_0_212 
* INOUT : br_0_212 
* INOUT : bl_0_213 
* INOUT : br_0_213 
* INOUT : bl_0_214 
* INOUT : br_0_214 
* INOUT : bl_0_215 
* INOUT : br_0_215 
* INOUT : bl_0_216 
* INOUT : br_0_216 
* INOUT : bl_0_217 
* INOUT : br_0_217 
* INOUT : bl_0_218 
* INOUT : br_0_218 
* INOUT : bl_0_219 
* INOUT : br_0_219 
* INOUT : bl_0_220 
* INOUT : br_0_220 
* INOUT : bl_0_221 
* INOUT : br_0_221 
* INOUT : bl_0_222 
* INOUT : br_0_222 
* INOUT : bl_0_223 
* INOUT : br_0_223 
* INOUT : bl_0_224 
* INOUT : br_0_224 
* INOUT : bl_0_225 
* INOUT : br_0_225 
* INOUT : bl_0_226 
* INOUT : br_0_226 
* INOUT : bl_0_227 
* INOUT : br_0_227 
* INOUT : bl_0_228 
* INOUT : br_0_228 
* INOUT : bl_0_229 
* INOUT : br_0_229 
* INOUT : bl_0_230 
* INOUT : br_0_230 
* INOUT : bl_0_231 
* INOUT : br_0_231 
* INOUT : bl_0_232 
* INOUT : br_0_232 
* INOUT : bl_0_233 
* INOUT : br_0_233 
* INOUT : bl_0_234 
* INOUT : br_0_234 
* INOUT : bl_0_235 
* INOUT : br_0_235 
* INOUT : bl_0_236 
* INOUT : br_0_236 
* INOUT : bl_0_237 
* INOUT : br_0_237 
* INOUT : bl_0_238 
* INOUT : br_0_238 
* INOUT : bl_0_239 
* INOUT : br_0_239 
* INOUT : bl_0_240 
* INOUT : br_0_240 
* INOUT : bl_0_241 
* INOUT : br_0_241 
* INOUT : bl_0_242 
* INOUT : br_0_242 
* INOUT : bl_0_243 
* INOUT : br_0_243 
* INOUT : bl_0_244 
* INOUT : br_0_244 
* INOUT : bl_0_245 
* INOUT : br_0_245 
* INOUT : bl_0_246 
* INOUT : br_0_246 
* INOUT : bl_0_247 
* INOUT : br_0_247 
* INOUT : bl_0_248 
* INOUT : br_0_248 
* INOUT : bl_0_249 
* INOUT : br_0_249 
* INOUT : bl_0_250 
* INOUT : br_0_250 
* INOUT : bl_0_251 
* INOUT : br_0_251 
* INOUT : bl_0_252 
* INOUT : br_0_252 
* INOUT : bl_0_253 
* INOUT : br_0_253 
* INOUT : bl_0_254 
* INOUT : br_0_254 
* INOUT : bl_0_255 
* INOUT : br_0_255 
* INOUT : bl_0_256 
* INOUT : br_0_256 
* INPUT : wl_0_0 
* POWER : vdd 
* GROUND: gnd 
Xbit_r0_c0
+ bl_0_0 br_0_0 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c1
+ bl_0_1 br_0_1 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c2
+ bl_0_2 br_0_2 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c3
+ bl_0_3 br_0_3 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c4
+ bl_0_4 br_0_4 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c5
+ bl_0_5 br_0_5 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c6
+ bl_0_6 br_0_6 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c7
+ bl_0_7 br_0_7 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c8
+ bl_0_8 br_0_8 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c9
+ bl_0_9 br_0_9 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c10
+ bl_0_10 br_0_10 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c11
+ bl_0_11 br_0_11 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c12
+ bl_0_12 br_0_12 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c13
+ bl_0_13 br_0_13 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c14
+ bl_0_14 br_0_14 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c15
+ bl_0_15 br_0_15 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c16
+ bl_0_16 br_0_16 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c17
+ bl_0_17 br_0_17 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c18
+ bl_0_18 br_0_18 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c19
+ bl_0_19 br_0_19 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c20
+ bl_0_20 br_0_20 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c21
+ bl_0_21 br_0_21 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c22
+ bl_0_22 br_0_22 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c23
+ bl_0_23 br_0_23 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c24
+ bl_0_24 br_0_24 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c25
+ bl_0_25 br_0_25 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c26
+ bl_0_26 br_0_26 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c27
+ bl_0_27 br_0_27 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c28
+ bl_0_28 br_0_28 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c29
+ bl_0_29 br_0_29 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c30
+ bl_0_30 br_0_30 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c31
+ bl_0_31 br_0_31 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c32
+ bl_0_32 br_0_32 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c33
+ bl_0_33 br_0_33 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c34
+ bl_0_34 br_0_34 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c35
+ bl_0_35 br_0_35 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c36
+ bl_0_36 br_0_36 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c37
+ bl_0_37 br_0_37 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c38
+ bl_0_38 br_0_38 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c39
+ bl_0_39 br_0_39 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c40
+ bl_0_40 br_0_40 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c41
+ bl_0_41 br_0_41 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c42
+ bl_0_42 br_0_42 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c43
+ bl_0_43 br_0_43 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c44
+ bl_0_44 br_0_44 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c45
+ bl_0_45 br_0_45 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c46
+ bl_0_46 br_0_46 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c47
+ bl_0_47 br_0_47 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c48
+ bl_0_48 br_0_48 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c49
+ bl_0_49 br_0_49 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c50
+ bl_0_50 br_0_50 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c51
+ bl_0_51 br_0_51 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c52
+ bl_0_52 br_0_52 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c53
+ bl_0_53 br_0_53 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c54
+ bl_0_54 br_0_54 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c55
+ bl_0_55 br_0_55 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c56
+ bl_0_56 br_0_56 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c57
+ bl_0_57 br_0_57 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c58
+ bl_0_58 br_0_58 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c59
+ bl_0_59 br_0_59 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c60
+ bl_0_60 br_0_60 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c61
+ bl_0_61 br_0_61 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c62
+ bl_0_62 br_0_62 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c63
+ bl_0_63 br_0_63 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c64
+ bl_0_64 br_0_64 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c65
+ bl_0_65 br_0_65 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c66
+ bl_0_66 br_0_66 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c67
+ bl_0_67 br_0_67 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c68
+ bl_0_68 br_0_68 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c69
+ bl_0_69 br_0_69 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c70
+ bl_0_70 br_0_70 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c71
+ bl_0_71 br_0_71 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c72
+ bl_0_72 br_0_72 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c73
+ bl_0_73 br_0_73 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c74
+ bl_0_74 br_0_74 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c75
+ bl_0_75 br_0_75 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c76
+ bl_0_76 br_0_76 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c77
+ bl_0_77 br_0_77 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c78
+ bl_0_78 br_0_78 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c79
+ bl_0_79 br_0_79 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c80
+ bl_0_80 br_0_80 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c81
+ bl_0_81 br_0_81 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c82
+ bl_0_82 br_0_82 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c83
+ bl_0_83 br_0_83 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c84
+ bl_0_84 br_0_84 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c85
+ bl_0_85 br_0_85 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c86
+ bl_0_86 br_0_86 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c87
+ bl_0_87 br_0_87 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c88
+ bl_0_88 br_0_88 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c89
+ bl_0_89 br_0_89 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c90
+ bl_0_90 br_0_90 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c91
+ bl_0_91 br_0_91 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c92
+ bl_0_92 br_0_92 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c93
+ bl_0_93 br_0_93 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c94
+ bl_0_94 br_0_94 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c95
+ bl_0_95 br_0_95 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c96
+ bl_0_96 br_0_96 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c97
+ bl_0_97 br_0_97 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c98
+ bl_0_98 br_0_98 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c99
+ bl_0_99 br_0_99 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c100
+ bl_0_100 br_0_100 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c101
+ bl_0_101 br_0_101 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c102
+ bl_0_102 br_0_102 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c103
+ bl_0_103 br_0_103 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c104
+ bl_0_104 br_0_104 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c105
+ bl_0_105 br_0_105 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c106
+ bl_0_106 br_0_106 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c107
+ bl_0_107 br_0_107 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c108
+ bl_0_108 br_0_108 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c109
+ bl_0_109 br_0_109 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c110
+ bl_0_110 br_0_110 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c111
+ bl_0_111 br_0_111 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c112
+ bl_0_112 br_0_112 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c113
+ bl_0_113 br_0_113 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c114
+ bl_0_114 br_0_114 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c115
+ bl_0_115 br_0_115 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c116
+ bl_0_116 br_0_116 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c117
+ bl_0_117 br_0_117 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c118
+ bl_0_118 br_0_118 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c119
+ bl_0_119 br_0_119 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c120
+ bl_0_120 br_0_120 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c121
+ bl_0_121 br_0_121 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c122
+ bl_0_122 br_0_122 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c123
+ bl_0_123 br_0_123 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c124
+ bl_0_124 br_0_124 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c125
+ bl_0_125 br_0_125 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c126
+ bl_0_126 br_0_126 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c127
+ bl_0_127 br_0_127 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c128
+ bl_0_128 br_0_128 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c129
+ bl_0_129 br_0_129 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c130
+ bl_0_130 br_0_130 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c131
+ bl_0_131 br_0_131 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c132
+ bl_0_132 br_0_132 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c133
+ bl_0_133 br_0_133 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c134
+ bl_0_134 br_0_134 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c135
+ bl_0_135 br_0_135 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c136
+ bl_0_136 br_0_136 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c137
+ bl_0_137 br_0_137 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c138
+ bl_0_138 br_0_138 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c139
+ bl_0_139 br_0_139 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c140
+ bl_0_140 br_0_140 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c141
+ bl_0_141 br_0_141 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c142
+ bl_0_142 br_0_142 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c143
+ bl_0_143 br_0_143 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c144
+ bl_0_144 br_0_144 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c145
+ bl_0_145 br_0_145 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c146
+ bl_0_146 br_0_146 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c147
+ bl_0_147 br_0_147 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c148
+ bl_0_148 br_0_148 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c149
+ bl_0_149 br_0_149 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c150
+ bl_0_150 br_0_150 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c151
+ bl_0_151 br_0_151 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c152
+ bl_0_152 br_0_152 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c153
+ bl_0_153 br_0_153 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c154
+ bl_0_154 br_0_154 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c155
+ bl_0_155 br_0_155 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c156
+ bl_0_156 br_0_156 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c157
+ bl_0_157 br_0_157 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c158
+ bl_0_158 br_0_158 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c159
+ bl_0_159 br_0_159 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c160
+ bl_0_160 br_0_160 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c161
+ bl_0_161 br_0_161 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c162
+ bl_0_162 br_0_162 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c163
+ bl_0_163 br_0_163 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c164
+ bl_0_164 br_0_164 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c165
+ bl_0_165 br_0_165 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c166
+ bl_0_166 br_0_166 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c167
+ bl_0_167 br_0_167 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c168
+ bl_0_168 br_0_168 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c169
+ bl_0_169 br_0_169 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c170
+ bl_0_170 br_0_170 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c171
+ bl_0_171 br_0_171 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c172
+ bl_0_172 br_0_172 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c173
+ bl_0_173 br_0_173 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c174
+ bl_0_174 br_0_174 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c175
+ bl_0_175 br_0_175 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c176
+ bl_0_176 br_0_176 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c177
+ bl_0_177 br_0_177 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c178
+ bl_0_178 br_0_178 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c179
+ bl_0_179 br_0_179 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c180
+ bl_0_180 br_0_180 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c181
+ bl_0_181 br_0_181 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c182
+ bl_0_182 br_0_182 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c183
+ bl_0_183 br_0_183 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c184
+ bl_0_184 br_0_184 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c185
+ bl_0_185 br_0_185 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c186
+ bl_0_186 br_0_186 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c187
+ bl_0_187 br_0_187 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c188
+ bl_0_188 br_0_188 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c189
+ bl_0_189 br_0_189 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c190
+ bl_0_190 br_0_190 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c191
+ bl_0_191 br_0_191 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c192
+ bl_0_192 br_0_192 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c193
+ bl_0_193 br_0_193 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c194
+ bl_0_194 br_0_194 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c195
+ bl_0_195 br_0_195 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c196
+ bl_0_196 br_0_196 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c197
+ bl_0_197 br_0_197 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c198
+ bl_0_198 br_0_198 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c199
+ bl_0_199 br_0_199 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c200
+ bl_0_200 br_0_200 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c201
+ bl_0_201 br_0_201 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c202
+ bl_0_202 br_0_202 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c203
+ bl_0_203 br_0_203 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c204
+ bl_0_204 br_0_204 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c205
+ bl_0_205 br_0_205 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c206
+ bl_0_206 br_0_206 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c207
+ bl_0_207 br_0_207 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c208
+ bl_0_208 br_0_208 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c209
+ bl_0_209 br_0_209 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c210
+ bl_0_210 br_0_210 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c211
+ bl_0_211 br_0_211 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c212
+ bl_0_212 br_0_212 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c213
+ bl_0_213 br_0_213 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c214
+ bl_0_214 br_0_214 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c215
+ bl_0_215 br_0_215 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c216
+ bl_0_216 br_0_216 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c217
+ bl_0_217 br_0_217 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c218
+ bl_0_218 br_0_218 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c219
+ bl_0_219 br_0_219 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c220
+ bl_0_220 br_0_220 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c221
+ bl_0_221 br_0_221 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c222
+ bl_0_222 br_0_222 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c223
+ bl_0_223 br_0_223 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c224
+ bl_0_224 br_0_224 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c225
+ bl_0_225 br_0_225 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c226
+ bl_0_226 br_0_226 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c227
+ bl_0_227 br_0_227 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c228
+ bl_0_228 br_0_228 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c229
+ bl_0_229 br_0_229 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c230
+ bl_0_230 br_0_230 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c231
+ bl_0_231 br_0_231 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c232
+ bl_0_232 br_0_232 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c233
+ bl_0_233 br_0_233 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c234
+ bl_0_234 br_0_234 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c235
+ bl_0_235 br_0_235 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c236
+ bl_0_236 br_0_236 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c237
+ bl_0_237 br_0_237 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c238
+ bl_0_238 br_0_238 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c239
+ bl_0_239 br_0_239 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c240
+ bl_0_240 br_0_240 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c241
+ bl_0_241 br_0_241 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c242
+ bl_0_242 br_0_242 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c243
+ bl_0_243 br_0_243 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c244
+ bl_0_244 br_0_244 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c245
+ bl_0_245 br_0_245 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c246
+ bl_0_246 br_0_246 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c247
+ bl_0_247 br_0_247 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c248
+ bl_0_248 br_0_248 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c249
+ bl_0_249 br_0_249 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c250
+ bl_0_250 br_0_250 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c251
+ bl_0_251 br_0_251 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c252
+ bl_0_252 br_0_252 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c253
+ bl_0_253 br_0_253 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c254
+ bl_0_254 br_0_254 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c255
+ bl_0_255 br_0_255 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c256
+ bl_0_256 br_0_256 wl_0_0 vdd gnd
+ dummy_cell_1rw
.ENDS sram_1rw0r0w_32_1024_freepdk45_dummy_array_0

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_dummy_array_3
+ bl_0_0 br_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7
+ wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16
+ wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24
+ wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32
+ wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40
+ wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48
+ wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56
+ wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64
+ wl_0_65 wl_0_66 wl_0_67 wl_0_68 wl_0_69 wl_0_70 wl_0_71 wl_0_72
+ wl_0_73 wl_0_74 wl_0_75 wl_0_76 wl_0_77 wl_0_78 wl_0_79 wl_0_80
+ wl_0_81 wl_0_82 wl_0_83 wl_0_84 wl_0_85 wl_0_86 wl_0_87 wl_0_88
+ wl_0_89 wl_0_90 wl_0_91 wl_0_92 wl_0_93 wl_0_94 wl_0_95 wl_0_96
+ wl_0_97 wl_0_98 wl_0_99 wl_0_100 wl_0_101 wl_0_102 wl_0_103 wl_0_104
+ wl_0_105 wl_0_106 wl_0_107 wl_0_108 wl_0_109 wl_0_110 wl_0_111
+ wl_0_112 wl_0_113 wl_0_114 wl_0_115 wl_0_116 wl_0_117 wl_0_118
+ wl_0_119 wl_0_120 wl_0_121 wl_0_122 wl_0_123 wl_0_124 wl_0_125
+ wl_0_126 wl_0_127 wl_0_128 wl_0_129 wl_0_130 vdd gnd
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* INPUT : wl_0_33 
* INPUT : wl_0_34 
* INPUT : wl_0_35 
* INPUT : wl_0_36 
* INPUT : wl_0_37 
* INPUT : wl_0_38 
* INPUT : wl_0_39 
* INPUT : wl_0_40 
* INPUT : wl_0_41 
* INPUT : wl_0_42 
* INPUT : wl_0_43 
* INPUT : wl_0_44 
* INPUT : wl_0_45 
* INPUT : wl_0_46 
* INPUT : wl_0_47 
* INPUT : wl_0_48 
* INPUT : wl_0_49 
* INPUT : wl_0_50 
* INPUT : wl_0_51 
* INPUT : wl_0_52 
* INPUT : wl_0_53 
* INPUT : wl_0_54 
* INPUT : wl_0_55 
* INPUT : wl_0_56 
* INPUT : wl_0_57 
* INPUT : wl_0_58 
* INPUT : wl_0_59 
* INPUT : wl_0_60 
* INPUT : wl_0_61 
* INPUT : wl_0_62 
* INPUT : wl_0_63 
* INPUT : wl_0_64 
* INPUT : wl_0_65 
* INPUT : wl_0_66 
* INPUT : wl_0_67 
* INPUT : wl_0_68 
* INPUT : wl_0_69 
* INPUT : wl_0_70 
* INPUT : wl_0_71 
* INPUT : wl_0_72 
* INPUT : wl_0_73 
* INPUT : wl_0_74 
* INPUT : wl_0_75 
* INPUT : wl_0_76 
* INPUT : wl_0_77 
* INPUT : wl_0_78 
* INPUT : wl_0_79 
* INPUT : wl_0_80 
* INPUT : wl_0_81 
* INPUT : wl_0_82 
* INPUT : wl_0_83 
* INPUT : wl_0_84 
* INPUT : wl_0_85 
* INPUT : wl_0_86 
* INPUT : wl_0_87 
* INPUT : wl_0_88 
* INPUT : wl_0_89 
* INPUT : wl_0_90 
* INPUT : wl_0_91 
* INPUT : wl_0_92 
* INPUT : wl_0_93 
* INPUT : wl_0_94 
* INPUT : wl_0_95 
* INPUT : wl_0_96 
* INPUT : wl_0_97 
* INPUT : wl_0_98 
* INPUT : wl_0_99 
* INPUT : wl_0_100 
* INPUT : wl_0_101 
* INPUT : wl_0_102 
* INPUT : wl_0_103 
* INPUT : wl_0_104 
* INPUT : wl_0_105 
* INPUT : wl_0_106 
* INPUT : wl_0_107 
* INPUT : wl_0_108 
* INPUT : wl_0_109 
* INPUT : wl_0_110 
* INPUT : wl_0_111 
* INPUT : wl_0_112 
* INPUT : wl_0_113 
* INPUT : wl_0_114 
* INPUT : wl_0_115 
* INPUT : wl_0_116 
* INPUT : wl_0_117 
* INPUT : wl_0_118 
* INPUT : wl_0_119 
* INPUT : wl_0_120 
* INPUT : wl_0_121 
* INPUT : wl_0_122 
* INPUT : wl_0_123 
* INPUT : wl_0_124 
* INPUT : wl_0_125 
* INPUT : wl_0_126 
* INPUT : wl_0_127 
* INPUT : wl_0_128 
* INPUT : wl_0_129 
* INPUT : wl_0_130 
* POWER : vdd 
* GROUND: gnd 
Xbit_r0_c0
+ bl_0_0 br_0_0 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r1_c0
+ bl_0_0 br_0_0 wl_0_1 vdd gnd
+ dummy_cell_1rw
Xbit_r2_c0
+ bl_0_0 br_0_0 wl_0_2 vdd gnd
+ dummy_cell_1rw
Xbit_r3_c0
+ bl_0_0 br_0_0 wl_0_3 vdd gnd
+ dummy_cell_1rw
Xbit_r4_c0
+ bl_0_0 br_0_0 wl_0_4 vdd gnd
+ dummy_cell_1rw
Xbit_r5_c0
+ bl_0_0 br_0_0 wl_0_5 vdd gnd
+ dummy_cell_1rw
Xbit_r6_c0
+ bl_0_0 br_0_0 wl_0_6 vdd gnd
+ dummy_cell_1rw
Xbit_r7_c0
+ bl_0_0 br_0_0 wl_0_7 vdd gnd
+ dummy_cell_1rw
Xbit_r8_c0
+ bl_0_0 br_0_0 wl_0_8 vdd gnd
+ dummy_cell_1rw
Xbit_r9_c0
+ bl_0_0 br_0_0 wl_0_9 vdd gnd
+ dummy_cell_1rw
Xbit_r10_c0
+ bl_0_0 br_0_0 wl_0_10 vdd gnd
+ dummy_cell_1rw
Xbit_r11_c0
+ bl_0_0 br_0_0 wl_0_11 vdd gnd
+ dummy_cell_1rw
Xbit_r12_c0
+ bl_0_0 br_0_0 wl_0_12 vdd gnd
+ dummy_cell_1rw
Xbit_r13_c0
+ bl_0_0 br_0_0 wl_0_13 vdd gnd
+ dummy_cell_1rw
Xbit_r14_c0
+ bl_0_0 br_0_0 wl_0_14 vdd gnd
+ dummy_cell_1rw
Xbit_r15_c0
+ bl_0_0 br_0_0 wl_0_15 vdd gnd
+ dummy_cell_1rw
Xbit_r16_c0
+ bl_0_0 br_0_0 wl_0_16 vdd gnd
+ dummy_cell_1rw
Xbit_r17_c0
+ bl_0_0 br_0_0 wl_0_17 vdd gnd
+ dummy_cell_1rw
Xbit_r18_c0
+ bl_0_0 br_0_0 wl_0_18 vdd gnd
+ dummy_cell_1rw
Xbit_r19_c0
+ bl_0_0 br_0_0 wl_0_19 vdd gnd
+ dummy_cell_1rw
Xbit_r20_c0
+ bl_0_0 br_0_0 wl_0_20 vdd gnd
+ dummy_cell_1rw
Xbit_r21_c0
+ bl_0_0 br_0_0 wl_0_21 vdd gnd
+ dummy_cell_1rw
Xbit_r22_c0
+ bl_0_0 br_0_0 wl_0_22 vdd gnd
+ dummy_cell_1rw
Xbit_r23_c0
+ bl_0_0 br_0_0 wl_0_23 vdd gnd
+ dummy_cell_1rw
Xbit_r24_c0
+ bl_0_0 br_0_0 wl_0_24 vdd gnd
+ dummy_cell_1rw
Xbit_r25_c0
+ bl_0_0 br_0_0 wl_0_25 vdd gnd
+ dummy_cell_1rw
Xbit_r26_c0
+ bl_0_0 br_0_0 wl_0_26 vdd gnd
+ dummy_cell_1rw
Xbit_r27_c0
+ bl_0_0 br_0_0 wl_0_27 vdd gnd
+ dummy_cell_1rw
Xbit_r28_c0
+ bl_0_0 br_0_0 wl_0_28 vdd gnd
+ dummy_cell_1rw
Xbit_r29_c0
+ bl_0_0 br_0_0 wl_0_29 vdd gnd
+ dummy_cell_1rw
Xbit_r30_c0
+ bl_0_0 br_0_0 wl_0_30 vdd gnd
+ dummy_cell_1rw
Xbit_r31_c0
+ bl_0_0 br_0_0 wl_0_31 vdd gnd
+ dummy_cell_1rw
Xbit_r32_c0
+ bl_0_0 br_0_0 wl_0_32 vdd gnd
+ dummy_cell_1rw
Xbit_r33_c0
+ bl_0_0 br_0_0 wl_0_33 vdd gnd
+ dummy_cell_1rw
Xbit_r34_c0
+ bl_0_0 br_0_0 wl_0_34 vdd gnd
+ dummy_cell_1rw
Xbit_r35_c0
+ bl_0_0 br_0_0 wl_0_35 vdd gnd
+ dummy_cell_1rw
Xbit_r36_c0
+ bl_0_0 br_0_0 wl_0_36 vdd gnd
+ dummy_cell_1rw
Xbit_r37_c0
+ bl_0_0 br_0_0 wl_0_37 vdd gnd
+ dummy_cell_1rw
Xbit_r38_c0
+ bl_0_0 br_0_0 wl_0_38 vdd gnd
+ dummy_cell_1rw
Xbit_r39_c0
+ bl_0_0 br_0_0 wl_0_39 vdd gnd
+ dummy_cell_1rw
Xbit_r40_c0
+ bl_0_0 br_0_0 wl_0_40 vdd gnd
+ dummy_cell_1rw
Xbit_r41_c0
+ bl_0_0 br_0_0 wl_0_41 vdd gnd
+ dummy_cell_1rw
Xbit_r42_c0
+ bl_0_0 br_0_0 wl_0_42 vdd gnd
+ dummy_cell_1rw
Xbit_r43_c0
+ bl_0_0 br_0_0 wl_0_43 vdd gnd
+ dummy_cell_1rw
Xbit_r44_c0
+ bl_0_0 br_0_0 wl_0_44 vdd gnd
+ dummy_cell_1rw
Xbit_r45_c0
+ bl_0_0 br_0_0 wl_0_45 vdd gnd
+ dummy_cell_1rw
Xbit_r46_c0
+ bl_0_0 br_0_0 wl_0_46 vdd gnd
+ dummy_cell_1rw
Xbit_r47_c0
+ bl_0_0 br_0_0 wl_0_47 vdd gnd
+ dummy_cell_1rw
Xbit_r48_c0
+ bl_0_0 br_0_0 wl_0_48 vdd gnd
+ dummy_cell_1rw
Xbit_r49_c0
+ bl_0_0 br_0_0 wl_0_49 vdd gnd
+ dummy_cell_1rw
Xbit_r50_c0
+ bl_0_0 br_0_0 wl_0_50 vdd gnd
+ dummy_cell_1rw
Xbit_r51_c0
+ bl_0_0 br_0_0 wl_0_51 vdd gnd
+ dummy_cell_1rw
Xbit_r52_c0
+ bl_0_0 br_0_0 wl_0_52 vdd gnd
+ dummy_cell_1rw
Xbit_r53_c0
+ bl_0_0 br_0_0 wl_0_53 vdd gnd
+ dummy_cell_1rw
Xbit_r54_c0
+ bl_0_0 br_0_0 wl_0_54 vdd gnd
+ dummy_cell_1rw
Xbit_r55_c0
+ bl_0_0 br_0_0 wl_0_55 vdd gnd
+ dummy_cell_1rw
Xbit_r56_c0
+ bl_0_0 br_0_0 wl_0_56 vdd gnd
+ dummy_cell_1rw
Xbit_r57_c0
+ bl_0_0 br_0_0 wl_0_57 vdd gnd
+ dummy_cell_1rw
Xbit_r58_c0
+ bl_0_0 br_0_0 wl_0_58 vdd gnd
+ dummy_cell_1rw
Xbit_r59_c0
+ bl_0_0 br_0_0 wl_0_59 vdd gnd
+ dummy_cell_1rw
Xbit_r60_c0
+ bl_0_0 br_0_0 wl_0_60 vdd gnd
+ dummy_cell_1rw
Xbit_r61_c0
+ bl_0_0 br_0_0 wl_0_61 vdd gnd
+ dummy_cell_1rw
Xbit_r62_c0
+ bl_0_0 br_0_0 wl_0_62 vdd gnd
+ dummy_cell_1rw
Xbit_r63_c0
+ bl_0_0 br_0_0 wl_0_63 vdd gnd
+ dummy_cell_1rw
Xbit_r64_c0
+ bl_0_0 br_0_0 wl_0_64 vdd gnd
+ dummy_cell_1rw
Xbit_r65_c0
+ bl_0_0 br_0_0 wl_0_65 vdd gnd
+ dummy_cell_1rw
Xbit_r66_c0
+ bl_0_0 br_0_0 wl_0_66 vdd gnd
+ dummy_cell_1rw
Xbit_r67_c0
+ bl_0_0 br_0_0 wl_0_67 vdd gnd
+ dummy_cell_1rw
Xbit_r68_c0
+ bl_0_0 br_0_0 wl_0_68 vdd gnd
+ dummy_cell_1rw
Xbit_r69_c0
+ bl_0_0 br_0_0 wl_0_69 vdd gnd
+ dummy_cell_1rw
Xbit_r70_c0
+ bl_0_0 br_0_0 wl_0_70 vdd gnd
+ dummy_cell_1rw
Xbit_r71_c0
+ bl_0_0 br_0_0 wl_0_71 vdd gnd
+ dummy_cell_1rw
Xbit_r72_c0
+ bl_0_0 br_0_0 wl_0_72 vdd gnd
+ dummy_cell_1rw
Xbit_r73_c0
+ bl_0_0 br_0_0 wl_0_73 vdd gnd
+ dummy_cell_1rw
Xbit_r74_c0
+ bl_0_0 br_0_0 wl_0_74 vdd gnd
+ dummy_cell_1rw
Xbit_r75_c0
+ bl_0_0 br_0_0 wl_0_75 vdd gnd
+ dummy_cell_1rw
Xbit_r76_c0
+ bl_0_0 br_0_0 wl_0_76 vdd gnd
+ dummy_cell_1rw
Xbit_r77_c0
+ bl_0_0 br_0_0 wl_0_77 vdd gnd
+ dummy_cell_1rw
Xbit_r78_c0
+ bl_0_0 br_0_0 wl_0_78 vdd gnd
+ dummy_cell_1rw
Xbit_r79_c0
+ bl_0_0 br_0_0 wl_0_79 vdd gnd
+ dummy_cell_1rw
Xbit_r80_c0
+ bl_0_0 br_0_0 wl_0_80 vdd gnd
+ dummy_cell_1rw
Xbit_r81_c0
+ bl_0_0 br_0_0 wl_0_81 vdd gnd
+ dummy_cell_1rw
Xbit_r82_c0
+ bl_0_0 br_0_0 wl_0_82 vdd gnd
+ dummy_cell_1rw
Xbit_r83_c0
+ bl_0_0 br_0_0 wl_0_83 vdd gnd
+ dummy_cell_1rw
Xbit_r84_c0
+ bl_0_0 br_0_0 wl_0_84 vdd gnd
+ dummy_cell_1rw
Xbit_r85_c0
+ bl_0_0 br_0_0 wl_0_85 vdd gnd
+ dummy_cell_1rw
Xbit_r86_c0
+ bl_0_0 br_0_0 wl_0_86 vdd gnd
+ dummy_cell_1rw
Xbit_r87_c0
+ bl_0_0 br_0_0 wl_0_87 vdd gnd
+ dummy_cell_1rw
Xbit_r88_c0
+ bl_0_0 br_0_0 wl_0_88 vdd gnd
+ dummy_cell_1rw
Xbit_r89_c0
+ bl_0_0 br_0_0 wl_0_89 vdd gnd
+ dummy_cell_1rw
Xbit_r90_c0
+ bl_0_0 br_0_0 wl_0_90 vdd gnd
+ dummy_cell_1rw
Xbit_r91_c0
+ bl_0_0 br_0_0 wl_0_91 vdd gnd
+ dummy_cell_1rw
Xbit_r92_c0
+ bl_0_0 br_0_0 wl_0_92 vdd gnd
+ dummy_cell_1rw
Xbit_r93_c0
+ bl_0_0 br_0_0 wl_0_93 vdd gnd
+ dummy_cell_1rw
Xbit_r94_c0
+ bl_0_0 br_0_0 wl_0_94 vdd gnd
+ dummy_cell_1rw
Xbit_r95_c0
+ bl_0_0 br_0_0 wl_0_95 vdd gnd
+ dummy_cell_1rw
Xbit_r96_c0
+ bl_0_0 br_0_0 wl_0_96 vdd gnd
+ dummy_cell_1rw
Xbit_r97_c0
+ bl_0_0 br_0_0 wl_0_97 vdd gnd
+ dummy_cell_1rw
Xbit_r98_c0
+ bl_0_0 br_0_0 wl_0_98 vdd gnd
+ dummy_cell_1rw
Xbit_r99_c0
+ bl_0_0 br_0_0 wl_0_99 vdd gnd
+ dummy_cell_1rw
Xbit_r100_c0
+ bl_0_0 br_0_0 wl_0_100 vdd gnd
+ dummy_cell_1rw
Xbit_r101_c0
+ bl_0_0 br_0_0 wl_0_101 vdd gnd
+ dummy_cell_1rw
Xbit_r102_c0
+ bl_0_0 br_0_0 wl_0_102 vdd gnd
+ dummy_cell_1rw
Xbit_r103_c0
+ bl_0_0 br_0_0 wl_0_103 vdd gnd
+ dummy_cell_1rw
Xbit_r104_c0
+ bl_0_0 br_0_0 wl_0_104 vdd gnd
+ dummy_cell_1rw
Xbit_r105_c0
+ bl_0_0 br_0_0 wl_0_105 vdd gnd
+ dummy_cell_1rw
Xbit_r106_c0
+ bl_0_0 br_0_0 wl_0_106 vdd gnd
+ dummy_cell_1rw
Xbit_r107_c0
+ bl_0_0 br_0_0 wl_0_107 vdd gnd
+ dummy_cell_1rw
Xbit_r108_c0
+ bl_0_0 br_0_0 wl_0_108 vdd gnd
+ dummy_cell_1rw
Xbit_r109_c0
+ bl_0_0 br_0_0 wl_0_109 vdd gnd
+ dummy_cell_1rw
Xbit_r110_c0
+ bl_0_0 br_0_0 wl_0_110 vdd gnd
+ dummy_cell_1rw
Xbit_r111_c0
+ bl_0_0 br_0_0 wl_0_111 vdd gnd
+ dummy_cell_1rw
Xbit_r112_c0
+ bl_0_0 br_0_0 wl_0_112 vdd gnd
+ dummy_cell_1rw
Xbit_r113_c0
+ bl_0_0 br_0_0 wl_0_113 vdd gnd
+ dummy_cell_1rw
Xbit_r114_c0
+ bl_0_0 br_0_0 wl_0_114 vdd gnd
+ dummy_cell_1rw
Xbit_r115_c0
+ bl_0_0 br_0_0 wl_0_115 vdd gnd
+ dummy_cell_1rw
Xbit_r116_c0
+ bl_0_0 br_0_0 wl_0_116 vdd gnd
+ dummy_cell_1rw
Xbit_r117_c0
+ bl_0_0 br_0_0 wl_0_117 vdd gnd
+ dummy_cell_1rw
Xbit_r118_c0
+ bl_0_0 br_0_0 wl_0_118 vdd gnd
+ dummy_cell_1rw
Xbit_r119_c0
+ bl_0_0 br_0_0 wl_0_119 vdd gnd
+ dummy_cell_1rw
Xbit_r120_c0
+ bl_0_0 br_0_0 wl_0_120 vdd gnd
+ dummy_cell_1rw
Xbit_r121_c0
+ bl_0_0 br_0_0 wl_0_121 vdd gnd
+ dummy_cell_1rw
Xbit_r122_c0
+ bl_0_0 br_0_0 wl_0_122 vdd gnd
+ dummy_cell_1rw
Xbit_r123_c0
+ bl_0_0 br_0_0 wl_0_123 vdd gnd
+ dummy_cell_1rw
Xbit_r124_c0
+ bl_0_0 br_0_0 wl_0_124 vdd gnd
+ dummy_cell_1rw
Xbit_r125_c0
+ bl_0_0 br_0_0 wl_0_125 vdd gnd
+ dummy_cell_1rw
Xbit_r126_c0
+ bl_0_0 br_0_0 wl_0_126 vdd gnd
+ dummy_cell_1rw
Xbit_r127_c0
+ bl_0_0 br_0_0 wl_0_127 vdd gnd
+ dummy_cell_1rw
Xbit_r128_c0
+ bl_0_0 br_0_0 wl_0_128 vdd gnd
+ dummy_cell_1rw
Xbit_r129_c0
+ bl_0_0 br_0_0 wl_0_129 vdd gnd
+ dummy_cell_1rw
Xbit_r130_c0
+ bl_0_0 br_0_0 wl_0_130 vdd gnd
+ dummy_cell_1rw
.ENDS sram_1rw0r0w_32_1024_freepdk45_dummy_array_3

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_capped_replica_bitcell_array
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64
+ bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68
+ bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72
+ bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76
+ bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80
+ bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84
+ bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88
+ bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92
+ bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96
+ bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100
+ bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104
+ br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107
+ bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111
+ br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114
+ bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118
+ br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121
+ bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125
+ br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128
+ bl_0_129 br_0_129 bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132
+ br_0_132 bl_0_133 br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135
+ bl_0_136 br_0_136 bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139
+ br_0_139 bl_0_140 br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142
+ bl_0_143 br_0_143 bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146
+ br_0_146 bl_0_147 br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149
+ bl_0_150 br_0_150 bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153
+ br_0_153 bl_0_154 br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156
+ bl_0_157 br_0_157 bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160
+ br_0_160 bl_0_161 br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163
+ bl_0_164 br_0_164 bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167
+ br_0_167 bl_0_168 br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170
+ bl_0_171 br_0_171 bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174
+ br_0_174 bl_0_175 br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177
+ bl_0_178 br_0_178 bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181
+ br_0_181 bl_0_182 br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184
+ bl_0_185 br_0_185 bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188
+ br_0_188 bl_0_189 br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191
+ bl_0_192 br_0_192 bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195
+ br_0_195 bl_0_196 br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198
+ bl_0_199 br_0_199 bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202
+ br_0_202 bl_0_203 br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205
+ bl_0_206 br_0_206 bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209
+ br_0_209 bl_0_210 br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212
+ bl_0_213 br_0_213 bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216
+ br_0_216 bl_0_217 br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219
+ bl_0_220 br_0_220 bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223
+ br_0_223 bl_0_224 br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226
+ bl_0_227 br_0_227 bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230
+ br_0_230 bl_0_231 br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233
+ bl_0_234 br_0_234 bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237
+ br_0_237 bl_0_238 br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240
+ bl_0_241 br_0_241 bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244
+ br_0_244 bl_0_245 br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247
+ bl_0_248 br_0_248 bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251
+ br_0_251 bl_0_252 br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254
+ bl_0_255 br_0_255 rbl_wl_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5
+ wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14
+ wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22
+ wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30
+ wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38
+ wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46
+ wl_0_47 wl_0_48 wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54
+ wl_0_55 wl_0_56 wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62
+ wl_0_63 wl_0_64 wl_0_65 wl_0_66 wl_0_67 wl_0_68 wl_0_69 wl_0_70
+ wl_0_71 wl_0_72 wl_0_73 wl_0_74 wl_0_75 wl_0_76 wl_0_77 wl_0_78
+ wl_0_79 wl_0_80 wl_0_81 wl_0_82 wl_0_83 wl_0_84 wl_0_85 wl_0_86
+ wl_0_87 wl_0_88 wl_0_89 wl_0_90 wl_0_91 wl_0_92 wl_0_93 wl_0_94
+ wl_0_95 wl_0_96 wl_0_97 wl_0_98 wl_0_99 wl_0_100 wl_0_101 wl_0_102
+ wl_0_103 wl_0_104 wl_0_105 wl_0_106 wl_0_107 wl_0_108 wl_0_109
+ wl_0_110 wl_0_111 wl_0_112 wl_0_113 wl_0_114 wl_0_115 wl_0_116
+ wl_0_117 wl_0_118 wl_0_119 wl_0_120 wl_0_121 wl_0_122 wl_0_123
+ wl_0_124 wl_0_125 wl_0_126 wl_0_127 vdd gnd
* INOUT : rbl_bl_0_0 
* INOUT : rbl_br_0_0 
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INOUT : bl_0_64 
* INOUT : br_0_64 
* INOUT : bl_0_65 
* INOUT : br_0_65 
* INOUT : bl_0_66 
* INOUT : br_0_66 
* INOUT : bl_0_67 
* INOUT : br_0_67 
* INOUT : bl_0_68 
* INOUT : br_0_68 
* INOUT : bl_0_69 
* INOUT : br_0_69 
* INOUT : bl_0_70 
* INOUT : br_0_70 
* INOUT : bl_0_71 
* INOUT : br_0_71 
* INOUT : bl_0_72 
* INOUT : br_0_72 
* INOUT : bl_0_73 
* INOUT : br_0_73 
* INOUT : bl_0_74 
* INOUT : br_0_74 
* INOUT : bl_0_75 
* INOUT : br_0_75 
* INOUT : bl_0_76 
* INOUT : br_0_76 
* INOUT : bl_0_77 
* INOUT : br_0_77 
* INOUT : bl_0_78 
* INOUT : br_0_78 
* INOUT : bl_0_79 
* INOUT : br_0_79 
* INOUT : bl_0_80 
* INOUT : br_0_80 
* INOUT : bl_0_81 
* INOUT : br_0_81 
* INOUT : bl_0_82 
* INOUT : br_0_82 
* INOUT : bl_0_83 
* INOUT : br_0_83 
* INOUT : bl_0_84 
* INOUT : br_0_84 
* INOUT : bl_0_85 
* INOUT : br_0_85 
* INOUT : bl_0_86 
* INOUT : br_0_86 
* INOUT : bl_0_87 
* INOUT : br_0_87 
* INOUT : bl_0_88 
* INOUT : br_0_88 
* INOUT : bl_0_89 
* INOUT : br_0_89 
* INOUT : bl_0_90 
* INOUT : br_0_90 
* INOUT : bl_0_91 
* INOUT : br_0_91 
* INOUT : bl_0_92 
* INOUT : br_0_92 
* INOUT : bl_0_93 
* INOUT : br_0_93 
* INOUT : bl_0_94 
* INOUT : br_0_94 
* INOUT : bl_0_95 
* INOUT : br_0_95 
* INOUT : bl_0_96 
* INOUT : br_0_96 
* INOUT : bl_0_97 
* INOUT : br_0_97 
* INOUT : bl_0_98 
* INOUT : br_0_98 
* INOUT : bl_0_99 
* INOUT : br_0_99 
* INOUT : bl_0_100 
* INOUT : br_0_100 
* INOUT : bl_0_101 
* INOUT : br_0_101 
* INOUT : bl_0_102 
* INOUT : br_0_102 
* INOUT : bl_0_103 
* INOUT : br_0_103 
* INOUT : bl_0_104 
* INOUT : br_0_104 
* INOUT : bl_0_105 
* INOUT : br_0_105 
* INOUT : bl_0_106 
* INOUT : br_0_106 
* INOUT : bl_0_107 
* INOUT : br_0_107 
* INOUT : bl_0_108 
* INOUT : br_0_108 
* INOUT : bl_0_109 
* INOUT : br_0_109 
* INOUT : bl_0_110 
* INOUT : br_0_110 
* INOUT : bl_0_111 
* INOUT : br_0_111 
* INOUT : bl_0_112 
* INOUT : br_0_112 
* INOUT : bl_0_113 
* INOUT : br_0_113 
* INOUT : bl_0_114 
* INOUT : br_0_114 
* INOUT : bl_0_115 
* INOUT : br_0_115 
* INOUT : bl_0_116 
* INOUT : br_0_116 
* INOUT : bl_0_117 
* INOUT : br_0_117 
* INOUT : bl_0_118 
* INOUT : br_0_118 
* INOUT : bl_0_119 
* INOUT : br_0_119 
* INOUT : bl_0_120 
* INOUT : br_0_120 
* INOUT : bl_0_121 
* INOUT : br_0_121 
* INOUT : bl_0_122 
* INOUT : br_0_122 
* INOUT : bl_0_123 
* INOUT : br_0_123 
* INOUT : bl_0_124 
* INOUT : br_0_124 
* INOUT : bl_0_125 
* INOUT : br_0_125 
* INOUT : bl_0_126 
* INOUT : br_0_126 
* INOUT : bl_0_127 
* INOUT : br_0_127 
* INOUT : bl_0_128 
* INOUT : br_0_128 
* INOUT : bl_0_129 
* INOUT : br_0_129 
* INOUT : bl_0_130 
* INOUT : br_0_130 
* INOUT : bl_0_131 
* INOUT : br_0_131 
* INOUT : bl_0_132 
* INOUT : br_0_132 
* INOUT : bl_0_133 
* INOUT : br_0_133 
* INOUT : bl_0_134 
* INOUT : br_0_134 
* INOUT : bl_0_135 
* INOUT : br_0_135 
* INOUT : bl_0_136 
* INOUT : br_0_136 
* INOUT : bl_0_137 
* INOUT : br_0_137 
* INOUT : bl_0_138 
* INOUT : br_0_138 
* INOUT : bl_0_139 
* INOUT : br_0_139 
* INOUT : bl_0_140 
* INOUT : br_0_140 
* INOUT : bl_0_141 
* INOUT : br_0_141 
* INOUT : bl_0_142 
* INOUT : br_0_142 
* INOUT : bl_0_143 
* INOUT : br_0_143 
* INOUT : bl_0_144 
* INOUT : br_0_144 
* INOUT : bl_0_145 
* INOUT : br_0_145 
* INOUT : bl_0_146 
* INOUT : br_0_146 
* INOUT : bl_0_147 
* INOUT : br_0_147 
* INOUT : bl_0_148 
* INOUT : br_0_148 
* INOUT : bl_0_149 
* INOUT : br_0_149 
* INOUT : bl_0_150 
* INOUT : br_0_150 
* INOUT : bl_0_151 
* INOUT : br_0_151 
* INOUT : bl_0_152 
* INOUT : br_0_152 
* INOUT : bl_0_153 
* INOUT : br_0_153 
* INOUT : bl_0_154 
* INOUT : br_0_154 
* INOUT : bl_0_155 
* INOUT : br_0_155 
* INOUT : bl_0_156 
* INOUT : br_0_156 
* INOUT : bl_0_157 
* INOUT : br_0_157 
* INOUT : bl_0_158 
* INOUT : br_0_158 
* INOUT : bl_0_159 
* INOUT : br_0_159 
* INOUT : bl_0_160 
* INOUT : br_0_160 
* INOUT : bl_0_161 
* INOUT : br_0_161 
* INOUT : bl_0_162 
* INOUT : br_0_162 
* INOUT : bl_0_163 
* INOUT : br_0_163 
* INOUT : bl_0_164 
* INOUT : br_0_164 
* INOUT : bl_0_165 
* INOUT : br_0_165 
* INOUT : bl_0_166 
* INOUT : br_0_166 
* INOUT : bl_0_167 
* INOUT : br_0_167 
* INOUT : bl_0_168 
* INOUT : br_0_168 
* INOUT : bl_0_169 
* INOUT : br_0_169 
* INOUT : bl_0_170 
* INOUT : br_0_170 
* INOUT : bl_0_171 
* INOUT : br_0_171 
* INOUT : bl_0_172 
* INOUT : br_0_172 
* INOUT : bl_0_173 
* INOUT : br_0_173 
* INOUT : bl_0_174 
* INOUT : br_0_174 
* INOUT : bl_0_175 
* INOUT : br_0_175 
* INOUT : bl_0_176 
* INOUT : br_0_176 
* INOUT : bl_0_177 
* INOUT : br_0_177 
* INOUT : bl_0_178 
* INOUT : br_0_178 
* INOUT : bl_0_179 
* INOUT : br_0_179 
* INOUT : bl_0_180 
* INOUT : br_0_180 
* INOUT : bl_0_181 
* INOUT : br_0_181 
* INOUT : bl_0_182 
* INOUT : br_0_182 
* INOUT : bl_0_183 
* INOUT : br_0_183 
* INOUT : bl_0_184 
* INOUT : br_0_184 
* INOUT : bl_0_185 
* INOUT : br_0_185 
* INOUT : bl_0_186 
* INOUT : br_0_186 
* INOUT : bl_0_187 
* INOUT : br_0_187 
* INOUT : bl_0_188 
* INOUT : br_0_188 
* INOUT : bl_0_189 
* INOUT : br_0_189 
* INOUT : bl_0_190 
* INOUT : br_0_190 
* INOUT : bl_0_191 
* INOUT : br_0_191 
* INOUT : bl_0_192 
* INOUT : br_0_192 
* INOUT : bl_0_193 
* INOUT : br_0_193 
* INOUT : bl_0_194 
* INOUT : br_0_194 
* INOUT : bl_0_195 
* INOUT : br_0_195 
* INOUT : bl_0_196 
* INOUT : br_0_196 
* INOUT : bl_0_197 
* INOUT : br_0_197 
* INOUT : bl_0_198 
* INOUT : br_0_198 
* INOUT : bl_0_199 
* INOUT : br_0_199 
* INOUT : bl_0_200 
* INOUT : br_0_200 
* INOUT : bl_0_201 
* INOUT : br_0_201 
* INOUT : bl_0_202 
* INOUT : br_0_202 
* INOUT : bl_0_203 
* INOUT : br_0_203 
* INOUT : bl_0_204 
* INOUT : br_0_204 
* INOUT : bl_0_205 
* INOUT : br_0_205 
* INOUT : bl_0_206 
* INOUT : br_0_206 
* INOUT : bl_0_207 
* INOUT : br_0_207 
* INOUT : bl_0_208 
* INOUT : br_0_208 
* INOUT : bl_0_209 
* INOUT : br_0_209 
* INOUT : bl_0_210 
* INOUT : br_0_210 
* INOUT : bl_0_211 
* INOUT : br_0_211 
* INOUT : bl_0_212 
* INOUT : br_0_212 
* INOUT : bl_0_213 
* INOUT : br_0_213 
* INOUT : bl_0_214 
* INOUT : br_0_214 
* INOUT : bl_0_215 
* INOUT : br_0_215 
* INOUT : bl_0_216 
* INOUT : br_0_216 
* INOUT : bl_0_217 
* INOUT : br_0_217 
* INOUT : bl_0_218 
* INOUT : br_0_218 
* INOUT : bl_0_219 
* INOUT : br_0_219 
* INOUT : bl_0_220 
* INOUT : br_0_220 
* INOUT : bl_0_221 
* INOUT : br_0_221 
* INOUT : bl_0_222 
* INOUT : br_0_222 
* INOUT : bl_0_223 
* INOUT : br_0_223 
* INOUT : bl_0_224 
* INOUT : br_0_224 
* INOUT : bl_0_225 
* INOUT : br_0_225 
* INOUT : bl_0_226 
* INOUT : br_0_226 
* INOUT : bl_0_227 
* INOUT : br_0_227 
* INOUT : bl_0_228 
* INOUT : br_0_228 
* INOUT : bl_0_229 
* INOUT : br_0_229 
* INOUT : bl_0_230 
* INOUT : br_0_230 
* INOUT : bl_0_231 
* INOUT : br_0_231 
* INOUT : bl_0_232 
* INOUT : br_0_232 
* INOUT : bl_0_233 
* INOUT : br_0_233 
* INOUT : bl_0_234 
* INOUT : br_0_234 
* INOUT : bl_0_235 
* INOUT : br_0_235 
* INOUT : bl_0_236 
* INOUT : br_0_236 
* INOUT : bl_0_237 
* INOUT : br_0_237 
* INOUT : bl_0_238 
* INOUT : br_0_238 
* INOUT : bl_0_239 
* INOUT : br_0_239 
* INOUT : bl_0_240 
* INOUT : br_0_240 
* INOUT : bl_0_241 
* INOUT : br_0_241 
* INOUT : bl_0_242 
* INOUT : br_0_242 
* INOUT : bl_0_243 
* INOUT : br_0_243 
* INOUT : bl_0_244 
* INOUT : br_0_244 
* INOUT : bl_0_245 
* INOUT : br_0_245 
* INOUT : bl_0_246 
* INOUT : br_0_246 
* INOUT : bl_0_247 
* INOUT : br_0_247 
* INOUT : bl_0_248 
* INOUT : br_0_248 
* INOUT : bl_0_249 
* INOUT : br_0_249 
* INOUT : bl_0_250 
* INOUT : br_0_250 
* INOUT : bl_0_251 
* INOUT : br_0_251 
* INOUT : bl_0_252 
* INOUT : br_0_252 
* INOUT : bl_0_253 
* INOUT : br_0_253 
* INOUT : bl_0_254 
* INOUT : br_0_254 
* INOUT : bl_0_255 
* INOUT : br_0_255 
* INPUT : rbl_wl_0_0 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* INPUT : wl_0_33 
* INPUT : wl_0_34 
* INPUT : wl_0_35 
* INPUT : wl_0_36 
* INPUT : wl_0_37 
* INPUT : wl_0_38 
* INPUT : wl_0_39 
* INPUT : wl_0_40 
* INPUT : wl_0_41 
* INPUT : wl_0_42 
* INPUT : wl_0_43 
* INPUT : wl_0_44 
* INPUT : wl_0_45 
* INPUT : wl_0_46 
* INPUT : wl_0_47 
* INPUT : wl_0_48 
* INPUT : wl_0_49 
* INPUT : wl_0_50 
* INPUT : wl_0_51 
* INPUT : wl_0_52 
* INPUT : wl_0_53 
* INPUT : wl_0_54 
* INPUT : wl_0_55 
* INPUT : wl_0_56 
* INPUT : wl_0_57 
* INPUT : wl_0_58 
* INPUT : wl_0_59 
* INPUT : wl_0_60 
* INPUT : wl_0_61 
* INPUT : wl_0_62 
* INPUT : wl_0_63 
* INPUT : wl_0_64 
* INPUT : wl_0_65 
* INPUT : wl_0_66 
* INPUT : wl_0_67 
* INPUT : wl_0_68 
* INPUT : wl_0_69 
* INPUT : wl_0_70 
* INPUT : wl_0_71 
* INPUT : wl_0_72 
* INPUT : wl_0_73 
* INPUT : wl_0_74 
* INPUT : wl_0_75 
* INPUT : wl_0_76 
* INPUT : wl_0_77 
* INPUT : wl_0_78 
* INPUT : wl_0_79 
* INPUT : wl_0_80 
* INPUT : wl_0_81 
* INPUT : wl_0_82 
* INPUT : wl_0_83 
* INPUT : wl_0_84 
* INPUT : wl_0_85 
* INPUT : wl_0_86 
* INPUT : wl_0_87 
* INPUT : wl_0_88 
* INPUT : wl_0_89 
* INPUT : wl_0_90 
* INPUT : wl_0_91 
* INPUT : wl_0_92 
* INPUT : wl_0_93 
* INPUT : wl_0_94 
* INPUT : wl_0_95 
* INPUT : wl_0_96 
* INPUT : wl_0_97 
* INPUT : wl_0_98 
* INPUT : wl_0_99 
* INPUT : wl_0_100 
* INPUT : wl_0_101 
* INPUT : wl_0_102 
* INPUT : wl_0_103 
* INPUT : wl_0_104 
* INPUT : wl_0_105 
* INPUT : wl_0_106 
* INPUT : wl_0_107 
* INPUT : wl_0_108 
* INPUT : wl_0_109 
* INPUT : wl_0_110 
* INPUT : wl_0_111 
* INPUT : wl_0_112 
* INPUT : wl_0_113 
* INPUT : wl_0_114 
* INPUT : wl_0_115 
* INPUT : wl_0_116 
* INPUT : wl_0_117 
* INPUT : wl_0_118 
* INPUT : wl_0_119 
* INPUT : wl_0_120 
* INPUT : wl_0_121 
* INPUT : wl_0_122 
* INPUT : wl_0_123 
* INPUT : wl_0_124 
* INPUT : wl_0_125 
* INPUT : wl_0_126 
* INPUT : wl_0_127 
* POWER : vdd 
* GROUND: gnd 
* rows: 128 cols: 256
* rbl: [1, 0] left_rbl: [0] right_rbl: []
Xreplica_bitcell_array
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64
+ bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68
+ bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72
+ bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76
+ bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80
+ bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84
+ bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88
+ bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92
+ bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96
+ bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100
+ bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104
+ br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107
+ bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111
+ br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114
+ bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118
+ br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121
+ bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125
+ br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128
+ bl_0_129 br_0_129 bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132
+ br_0_132 bl_0_133 br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135
+ bl_0_136 br_0_136 bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139
+ br_0_139 bl_0_140 br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142
+ bl_0_143 br_0_143 bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146
+ br_0_146 bl_0_147 br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149
+ bl_0_150 br_0_150 bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153
+ br_0_153 bl_0_154 br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156
+ bl_0_157 br_0_157 bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160
+ br_0_160 bl_0_161 br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163
+ bl_0_164 br_0_164 bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167
+ br_0_167 bl_0_168 br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170
+ bl_0_171 br_0_171 bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174
+ br_0_174 bl_0_175 br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177
+ bl_0_178 br_0_178 bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181
+ br_0_181 bl_0_182 br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184
+ bl_0_185 br_0_185 bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188
+ br_0_188 bl_0_189 br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191
+ bl_0_192 br_0_192 bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195
+ br_0_195 bl_0_196 br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198
+ bl_0_199 br_0_199 bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202
+ br_0_202 bl_0_203 br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205
+ bl_0_206 br_0_206 bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209
+ br_0_209 bl_0_210 br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212
+ bl_0_213 br_0_213 bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216
+ br_0_216 bl_0_217 br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219
+ bl_0_220 br_0_220 bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223
+ br_0_223 bl_0_224 br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226
+ bl_0_227 br_0_227 bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230
+ br_0_230 bl_0_231 br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233
+ bl_0_234 br_0_234 bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237
+ br_0_237 bl_0_238 br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240
+ bl_0_241 br_0_241 bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244
+ br_0_244 bl_0_245 br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247
+ bl_0_248 br_0_248 bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251
+ br_0_251 bl_0_252 br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254
+ bl_0_255 br_0_255 rbl_wl_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5
+ wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14
+ wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22
+ wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30
+ wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38
+ wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46
+ wl_0_47 wl_0_48 wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54
+ wl_0_55 wl_0_56 wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62
+ wl_0_63 wl_0_64 wl_0_65 wl_0_66 wl_0_67 wl_0_68 wl_0_69 wl_0_70
+ wl_0_71 wl_0_72 wl_0_73 wl_0_74 wl_0_75 wl_0_76 wl_0_77 wl_0_78
+ wl_0_79 wl_0_80 wl_0_81 wl_0_82 wl_0_83 wl_0_84 wl_0_85 wl_0_86
+ wl_0_87 wl_0_88 wl_0_89 wl_0_90 wl_0_91 wl_0_92 wl_0_93 wl_0_94
+ wl_0_95 wl_0_96 wl_0_97 wl_0_98 wl_0_99 wl_0_100 wl_0_101 wl_0_102
+ wl_0_103 wl_0_104 wl_0_105 wl_0_106 wl_0_107 wl_0_108 wl_0_109
+ wl_0_110 wl_0_111 wl_0_112 wl_0_113 wl_0_114 wl_0_115 wl_0_116
+ wl_0_117 wl_0_118 wl_0_119 wl_0_120 wl_0_121 wl_0_122 wl_0_123
+ wl_0_124 wl_0_125 wl_0_126 wl_0_127 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_replica_bitcell_array
Xdummy_row_bot
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64
+ bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68
+ bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72
+ bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76
+ bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80
+ bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84
+ bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88
+ bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92
+ bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96
+ bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100
+ bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104
+ br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107
+ bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111
+ br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114
+ bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118
+ br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121
+ bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125
+ br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128
+ bl_0_129 br_0_129 bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132
+ br_0_132 bl_0_133 br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135
+ bl_0_136 br_0_136 bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139
+ br_0_139 bl_0_140 br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142
+ bl_0_143 br_0_143 bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146
+ br_0_146 bl_0_147 br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149
+ bl_0_150 br_0_150 bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153
+ br_0_153 bl_0_154 br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156
+ bl_0_157 br_0_157 bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160
+ br_0_160 bl_0_161 br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163
+ bl_0_164 br_0_164 bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167
+ br_0_167 bl_0_168 br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170
+ bl_0_171 br_0_171 bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174
+ br_0_174 bl_0_175 br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177
+ bl_0_178 br_0_178 bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181
+ br_0_181 bl_0_182 br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184
+ bl_0_185 br_0_185 bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188
+ br_0_188 bl_0_189 br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191
+ bl_0_192 br_0_192 bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195
+ br_0_195 bl_0_196 br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198
+ bl_0_199 br_0_199 bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202
+ br_0_202 bl_0_203 br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205
+ bl_0_206 br_0_206 bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209
+ br_0_209 bl_0_210 br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212
+ bl_0_213 br_0_213 bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216
+ br_0_216 bl_0_217 br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219
+ bl_0_220 br_0_220 bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223
+ br_0_223 bl_0_224 br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226
+ bl_0_227 br_0_227 bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230
+ br_0_230 bl_0_231 br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233
+ bl_0_234 br_0_234 bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237
+ br_0_237 bl_0_238 br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240
+ bl_0_241 br_0_241 bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244
+ br_0_244 bl_0_245 br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247
+ bl_0_248 br_0_248 bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251
+ br_0_251 bl_0_252 br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254
+ bl_0_255 br_0_255 gnd vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_dummy_array_1
Xdummy_row_top
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64
+ bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68
+ bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72
+ bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76
+ bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80
+ bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84
+ bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88
+ bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92
+ bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96
+ bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100
+ bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104
+ br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107
+ bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111
+ br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114
+ bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118
+ br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121
+ bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125
+ br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128
+ bl_0_129 br_0_129 bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132
+ br_0_132 bl_0_133 br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135
+ bl_0_136 br_0_136 bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139
+ br_0_139 bl_0_140 br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142
+ bl_0_143 br_0_143 bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146
+ br_0_146 bl_0_147 br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149
+ bl_0_150 br_0_150 bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153
+ br_0_153 bl_0_154 br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156
+ bl_0_157 br_0_157 bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160
+ br_0_160 bl_0_161 br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163
+ bl_0_164 br_0_164 bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167
+ br_0_167 bl_0_168 br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170
+ bl_0_171 br_0_171 bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174
+ br_0_174 bl_0_175 br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177
+ bl_0_178 br_0_178 bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181
+ br_0_181 bl_0_182 br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184
+ bl_0_185 br_0_185 bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188
+ br_0_188 bl_0_189 br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191
+ bl_0_192 br_0_192 bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195
+ br_0_195 bl_0_196 br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198
+ bl_0_199 br_0_199 bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202
+ br_0_202 bl_0_203 br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205
+ bl_0_206 br_0_206 bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209
+ br_0_209 bl_0_210 br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212
+ bl_0_213 br_0_213 bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216
+ br_0_216 bl_0_217 br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219
+ bl_0_220 br_0_220 bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223
+ br_0_223 bl_0_224 br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226
+ bl_0_227 br_0_227 bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230
+ br_0_230 bl_0_231 br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233
+ bl_0_234 br_0_234 bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237
+ br_0_237 bl_0_238 br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240
+ bl_0_241 br_0_241 bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244
+ br_0_244 bl_0_245 br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247
+ bl_0_248 br_0_248 bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251
+ br_0_251 bl_0_252 br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254
+ bl_0_255 br_0_255 gnd vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_dummy_array_0
Xdummy_col_left
+ dummy_left_bl_0_0 dummy_left_br_0_0 gnd rbl_wl_0_0 wl_0_0 wl_0_1
+ wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10
+ wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18
+ wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26
+ wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34
+ wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42
+ wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50
+ wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57 wl_0_58
+ wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 wl_0_65 wl_0_66
+ wl_0_67 wl_0_68 wl_0_69 wl_0_70 wl_0_71 wl_0_72 wl_0_73 wl_0_74
+ wl_0_75 wl_0_76 wl_0_77 wl_0_78 wl_0_79 wl_0_80 wl_0_81 wl_0_82
+ wl_0_83 wl_0_84 wl_0_85 wl_0_86 wl_0_87 wl_0_88 wl_0_89 wl_0_90
+ wl_0_91 wl_0_92 wl_0_93 wl_0_94 wl_0_95 wl_0_96 wl_0_97 wl_0_98
+ wl_0_99 wl_0_100 wl_0_101 wl_0_102 wl_0_103 wl_0_104 wl_0_105 wl_0_106
+ wl_0_107 wl_0_108 wl_0_109 wl_0_110 wl_0_111 wl_0_112 wl_0_113
+ wl_0_114 wl_0_115 wl_0_116 wl_0_117 wl_0_118 wl_0_119 wl_0_120
+ wl_0_121 wl_0_122 wl_0_123 wl_0_124 wl_0_125 wl_0_126 wl_0_127 gnd vdd
+ gnd
+ sram_1rw0r0w_32_1024_freepdk45_dummy_array_2
Xdummy_col_right
+ dummy_right_bl_0_0 dummy_right_br_0_0 gnd rbl_wl_0_0 wl_0_0 wl_0_1
+ wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10
+ wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18
+ wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26
+ wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34
+ wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42
+ wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50
+ wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57 wl_0_58
+ wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 wl_0_65 wl_0_66
+ wl_0_67 wl_0_68 wl_0_69 wl_0_70 wl_0_71 wl_0_72 wl_0_73 wl_0_74
+ wl_0_75 wl_0_76 wl_0_77 wl_0_78 wl_0_79 wl_0_80 wl_0_81 wl_0_82
+ wl_0_83 wl_0_84 wl_0_85 wl_0_86 wl_0_87 wl_0_88 wl_0_89 wl_0_90
+ wl_0_91 wl_0_92 wl_0_93 wl_0_94 wl_0_95 wl_0_96 wl_0_97 wl_0_98
+ wl_0_99 wl_0_100 wl_0_101 wl_0_102 wl_0_103 wl_0_104 wl_0_105 wl_0_106
+ wl_0_107 wl_0_108 wl_0_109 wl_0_110 wl_0_111 wl_0_112 wl_0_113
+ wl_0_114 wl_0_115 wl_0_116 wl_0_117 wl_0_118 wl_0_119 wl_0_120
+ wl_0_121 wl_0_122 wl_0_123 wl_0_124 wl_0_125 wl_0_126 wl_0_127 gnd vdd
+ gnd
+ sram_1rw0r0w_32_1024_freepdk45_dummy_array_3
.ENDS sram_1rw0r0w_32_1024_freepdk45_capped_replica_bitcell_array

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_precharge_0
+ bl br en_bar vdd
* OUTPUT: bl 
* OUTPUT: br 
* INPUT : en_bar 
* POWER : vdd 
Mlower_pmos bl en_bar br vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mupper_pmos1 bl en_bar vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mupper_pmos2 br en_bar vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
.ENDS sram_1rw0r0w_32_1024_freepdk45_precharge_0

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_precharge_array
+ bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6
+ bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12
+ bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18
+ br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23
+ bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29
+ br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34
+ bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40
+ br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45
+ bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51
+ br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56
+ bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62
+ br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67
+ bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73
+ br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78
+ bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84
+ br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89
+ bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95
+ br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100
+ bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105
+ bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110
+ bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115
+ bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120
+ bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125
+ bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130
+ bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135
+ bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140
+ bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145
+ bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150
+ bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155
+ bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160
+ bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165
+ bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170
+ bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175
+ bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180
+ bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185
+ bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190
+ bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195
+ bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200
+ bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205
+ bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210
+ bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215
+ bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220
+ bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225
+ bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230
+ bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235
+ bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240
+ bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245
+ bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250
+ bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255
+ bl_256 br_256 en_bar vdd
* OUTPUT: bl_0 
* OUTPUT: br_0 
* OUTPUT: bl_1 
* OUTPUT: br_1 
* OUTPUT: bl_2 
* OUTPUT: br_2 
* OUTPUT: bl_3 
* OUTPUT: br_3 
* OUTPUT: bl_4 
* OUTPUT: br_4 
* OUTPUT: bl_5 
* OUTPUT: br_5 
* OUTPUT: bl_6 
* OUTPUT: br_6 
* OUTPUT: bl_7 
* OUTPUT: br_7 
* OUTPUT: bl_8 
* OUTPUT: br_8 
* OUTPUT: bl_9 
* OUTPUT: br_9 
* OUTPUT: bl_10 
* OUTPUT: br_10 
* OUTPUT: bl_11 
* OUTPUT: br_11 
* OUTPUT: bl_12 
* OUTPUT: br_12 
* OUTPUT: bl_13 
* OUTPUT: br_13 
* OUTPUT: bl_14 
* OUTPUT: br_14 
* OUTPUT: bl_15 
* OUTPUT: br_15 
* OUTPUT: bl_16 
* OUTPUT: br_16 
* OUTPUT: bl_17 
* OUTPUT: br_17 
* OUTPUT: bl_18 
* OUTPUT: br_18 
* OUTPUT: bl_19 
* OUTPUT: br_19 
* OUTPUT: bl_20 
* OUTPUT: br_20 
* OUTPUT: bl_21 
* OUTPUT: br_21 
* OUTPUT: bl_22 
* OUTPUT: br_22 
* OUTPUT: bl_23 
* OUTPUT: br_23 
* OUTPUT: bl_24 
* OUTPUT: br_24 
* OUTPUT: bl_25 
* OUTPUT: br_25 
* OUTPUT: bl_26 
* OUTPUT: br_26 
* OUTPUT: bl_27 
* OUTPUT: br_27 
* OUTPUT: bl_28 
* OUTPUT: br_28 
* OUTPUT: bl_29 
* OUTPUT: br_29 
* OUTPUT: bl_30 
* OUTPUT: br_30 
* OUTPUT: bl_31 
* OUTPUT: br_31 
* OUTPUT: bl_32 
* OUTPUT: br_32 
* OUTPUT: bl_33 
* OUTPUT: br_33 
* OUTPUT: bl_34 
* OUTPUT: br_34 
* OUTPUT: bl_35 
* OUTPUT: br_35 
* OUTPUT: bl_36 
* OUTPUT: br_36 
* OUTPUT: bl_37 
* OUTPUT: br_37 
* OUTPUT: bl_38 
* OUTPUT: br_38 
* OUTPUT: bl_39 
* OUTPUT: br_39 
* OUTPUT: bl_40 
* OUTPUT: br_40 
* OUTPUT: bl_41 
* OUTPUT: br_41 
* OUTPUT: bl_42 
* OUTPUT: br_42 
* OUTPUT: bl_43 
* OUTPUT: br_43 
* OUTPUT: bl_44 
* OUTPUT: br_44 
* OUTPUT: bl_45 
* OUTPUT: br_45 
* OUTPUT: bl_46 
* OUTPUT: br_46 
* OUTPUT: bl_47 
* OUTPUT: br_47 
* OUTPUT: bl_48 
* OUTPUT: br_48 
* OUTPUT: bl_49 
* OUTPUT: br_49 
* OUTPUT: bl_50 
* OUTPUT: br_50 
* OUTPUT: bl_51 
* OUTPUT: br_51 
* OUTPUT: bl_52 
* OUTPUT: br_52 
* OUTPUT: bl_53 
* OUTPUT: br_53 
* OUTPUT: bl_54 
* OUTPUT: br_54 
* OUTPUT: bl_55 
* OUTPUT: br_55 
* OUTPUT: bl_56 
* OUTPUT: br_56 
* OUTPUT: bl_57 
* OUTPUT: br_57 
* OUTPUT: bl_58 
* OUTPUT: br_58 
* OUTPUT: bl_59 
* OUTPUT: br_59 
* OUTPUT: bl_60 
* OUTPUT: br_60 
* OUTPUT: bl_61 
* OUTPUT: br_61 
* OUTPUT: bl_62 
* OUTPUT: br_62 
* OUTPUT: bl_63 
* OUTPUT: br_63 
* OUTPUT: bl_64 
* OUTPUT: br_64 
* OUTPUT: bl_65 
* OUTPUT: br_65 
* OUTPUT: bl_66 
* OUTPUT: br_66 
* OUTPUT: bl_67 
* OUTPUT: br_67 
* OUTPUT: bl_68 
* OUTPUT: br_68 
* OUTPUT: bl_69 
* OUTPUT: br_69 
* OUTPUT: bl_70 
* OUTPUT: br_70 
* OUTPUT: bl_71 
* OUTPUT: br_71 
* OUTPUT: bl_72 
* OUTPUT: br_72 
* OUTPUT: bl_73 
* OUTPUT: br_73 
* OUTPUT: bl_74 
* OUTPUT: br_74 
* OUTPUT: bl_75 
* OUTPUT: br_75 
* OUTPUT: bl_76 
* OUTPUT: br_76 
* OUTPUT: bl_77 
* OUTPUT: br_77 
* OUTPUT: bl_78 
* OUTPUT: br_78 
* OUTPUT: bl_79 
* OUTPUT: br_79 
* OUTPUT: bl_80 
* OUTPUT: br_80 
* OUTPUT: bl_81 
* OUTPUT: br_81 
* OUTPUT: bl_82 
* OUTPUT: br_82 
* OUTPUT: bl_83 
* OUTPUT: br_83 
* OUTPUT: bl_84 
* OUTPUT: br_84 
* OUTPUT: bl_85 
* OUTPUT: br_85 
* OUTPUT: bl_86 
* OUTPUT: br_86 
* OUTPUT: bl_87 
* OUTPUT: br_87 
* OUTPUT: bl_88 
* OUTPUT: br_88 
* OUTPUT: bl_89 
* OUTPUT: br_89 
* OUTPUT: bl_90 
* OUTPUT: br_90 
* OUTPUT: bl_91 
* OUTPUT: br_91 
* OUTPUT: bl_92 
* OUTPUT: br_92 
* OUTPUT: bl_93 
* OUTPUT: br_93 
* OUTPUT: bl_94 
* OUTPUT: br_94 
* OUTPUT: bl_95 
* OUTPUT: br_95 
* OUTPUT: bl_96 
* OUTPUT: br_96 
* OUTPUT: bl_97 
* OUTPUT: br_97 
* OUTPUT: bl_98 
* OUTPUT: br_98 
* OUTPUT: bl_99 
* OUTPUT: br_99 
* OUTPUT: bl_100 
* OUTPUT: br_100 
* OUTPUT: bl_101 
* OUTPUT: br_101 
* OUTPUT: bl_102 
* OUTPUT: br_102 
* OUTPUT: bl_103 
* OUTPUT: br_103 
* OUTPUT: bl_104 
* OUTPUT: br_104 
* OUTPUT: bl_105 
* OUTPUT: br_105 
* OUTPUT: bl_106 
* OUTPUT: br_106 
* OUTPUT: bl_107 
* OUTPUT: br_107 
* OUTPUT: bl_108 
* OUTPUT: br_108 
* OUTPUT: bl_109 
* OUTPUT: br_109 
* OUTPUT: bl_110 
* OUTPUT: br_110 
* OUTPUT: bl_111 
* OUTPUT: br_111 
* OUTPUT: bl_112 
* OUTPUT: br_112 
* OUTPUT: bl_113 
* OUTPUT: br_113 
* OUTPUT: bl_114 
* OUTPUT: br_114 
* OUTPUT: bl_115 
* OUTPUT: br_115 
* OUTPUT: bl_116 
* OUTPUT: br_116 
* OUTPUT: bl_117 
* OUTPUT: br_117 
* OUTPUT: bl_118 
* OUTPUT: br_118 
* OUTPUT: bl_119 
* OUTPUT: br_119 
* OUTPUT: bl_120 
* OUTPUT: br_120 
* OUTPUT: bl_121 
* OUTPUT: br_121 
* OUTPUT: bl_122 
* OUTPUT: br_122 
* OUTPUT: bl_123 
* OUTPUT: br_123 
* OUTPUT: bl_124 
* OUTPUT: br_124 
* OUTPUT: bl_125 
* OUTPUT: br_125 
* OUTPUT: bl_126 
* OUTPUT: br_126 
* OUTPUT: bl_127 
* OUTPUT: br_127 
* OUTPUT: bl_128 
* OUTPUT: br_128 
* OUTPUT: bl_129 
* OUTPUT: br_129 
* OUTPUT: bl_130 
* OUTPUT: br_130 
* OUTPUT: bl_131 
* OUTPUT: br_131 
* OUTPUT: bl_132 
* OUTPUT: br_132 
* OUTPUT: bl_133 
* OUTPUT: br_133 
* OUTPUT: bl_134 
* OUTPUT: br_134 
* OUTPUT: bl_135 
* OUTPUT: br_135 
* OUTPUT: bl_136 
* OUTPUT: br_136 
* OUTPUT: bl_137 
* OUTPUT: br_137 
* OUTPUT: bl_138 
* OUTPUT: br_138 
* OUTPUT: bl_139 
* OUTPUT: br_139 
* OUTPUT: bl_140 
* OUTPUT: br_140 
* OUTPUT: bl_141 
* OUTPUT: br_141 
* OUTPUT: bl_142 
* OUTPUT: br_142 
* OUTPUT: bl_143 
* OUTPUT: br_143 
* OUTPUT: bl_144 
* OUTPUT: br_144 
* OUTPUT: bl_145 
* OUTPUT: br_145 
* OUTPUT: bl_146 
* OUTPUT: br_146 
* OUTPUT: bl_147 
* OUTPUT: br_147 
* OUTPUT: bl_148 
* OUTPUT: br_148 
* OUTPUT: bl_149 
* OUTPUT: br_149 
* OUTPUT: bl_150 
* OUTPUT: br_150 
* OUTPUT: bl_151 
* OUTPUT: br_151 
* OUTPUT: bl_152 
* OUTPUT: br_152 
* OUTPUT: bl_153 
* OUTPUT: br_153 
* OUTPUT: bl_154 
* OUTPUT: br_154 
* OUTPUT: bl_155 
* OUTPUT: br_155 
* OUTPUT: bl_156 
* OUTPUT: br_156 
* OUTPUT: bl_157 
* OUTPUT: br_157 
* OUTPUT: bl_158 
* OUTPUT: br_158 
* OUTPUT: bl_159 
* OUTPUT: br_159 
* OUTPUT: bl_160 
* OUTPUT: br_160 
* OUTPUT: bl_161 
* OUTPUT: br_161 
* OUTPUT: bl_162 
* OUTPUT: br_162 
* OUTPUT: bl_163 
* OUTPUT: br_163 
* OUTPUT: bl_164 
* OUTPUT: br_164 
* OUTPUT: bl_165 
* OUTPUT: br_165 
* OUTPUT: bl_166 
* OUTPUT: br_166 
* OUTPUT: bl_167 
* OUTPUT: br_167 
* OUTPUT: bl_168 
* OUTPUT: br_168 
* OUTPUT: bl_169 
* OUTPUT: br_169 
* OUTPUT: bl_170 
* OUTPUT: br_170 
* OUTPUT: bl_171 
* OUTPUT: br_171 
* OUTPUT: bl_172 
* OUTPUT: br_172 
* OUTPUT: bl_173 
* OUTPUT: br_173 
* OUTPUT: bl_174 
* OUTPUT: br_174 
* OUTPUT: bl_175 
* OUTPUT: br_175 
* OUTPUT: bl_176 
* OUTPUT: br_176 
* OUTPUT: bl_177 
* OUTPUT: br_177 
* OUTPUT: bl_178 
* OUTPUT: br_178 
* OUTPUT: bl_179 
* OUTPUT: br_179 
* OUTPUT: bl_180 
* OUTPUT: br_180 
* OUTPUT: bl_181 
* OUTPUT: br_181 
* OUTPUT: bl_182 
* OUTPUT: br_182 
* OUTPUT: bl_183 
* OUTPUT: br_183 
* OUTPUT: bl_184 
* OUTPUT: br_184 
* OUTPUT: bl_185 
* OUTPUT: br_185 
* OUTPUT: bl_186 
* OUTPUT: br_186 
* OUTPUT: bl_187 
* OUTPUT: br_187 
* OUTPUT: bl_188 
* OUTPUT: br_188 
* OUTPUT: bl_189 
* OUTPUT: br_189 
* OUTPUT: bl_190 
* OUTPUT: br_190 
* OUTPUT: bl_191 
* OUTPUT: br_191 
* OUTPUT: bl_192 
* OUTPUT: br_192 
* OUTPUT: bl_193 
* OUTPUT: br_193 
* OUTPUT: bl_194 
* OUTPUT: br_194 
* OUTPUT: bl_195 
* OUTPUT: br_195 
* OUTPUT: bl_196 
* OUTPUT: br_196 
* OUTPUT: bl_197 
* OUTPUT: br_197 
* OUTPUT: bl_198 
* OUTPUT: br_198 
* OUTPUT: bl_199 
* OUTPUT: br_199 
* OUTPUT: bl_200 
* OUTPUT: br_200 
* OUTPUT: bl_201 
* OUTPUT: br_201 
* OUTPUT: bl_202 
* OUTPUT: br_202 
* OUTPUT: bl_203 
* OUTPUT: br_203 
* OUTPUT: bl_204 
* OUTPUT: br_204 
* OUTPUT: bl_205 
* OUTPUT: br_205 
* OUTPUT: bl_206 
* OUTPUT: br_206 
* OUTPUT: bl_207 
* OUTPUT: br_207 
* OUTPUT: bl_208 
* OUTPUT: br_208 
* OUTPUT: bl_209 
* OUTPUT: br_209 
* OUTPUT: bl_210 
* OUTPUT: br_210 
* OUTPUT: bl_211 
* OUTPUT: br_211 
* OUTPUT: bl_212 
* OUTPUT: br_212 
* OUTPUT: bl_213 
* OUTPUT: br_213 
* OUTPUT: bl_214 
* OUTPUT: br_214 
* OUTPUT: bl_215 
* OUTPUT: br_215 
* OUTPUT: bl_216 
* OUTPUT: br_216 
* OUTPUT: bl_217 
* OUTPUT: br_217 
* OUTPUT: bl_218 
* OUTPUT: br_218 
* OUTPUT: bl_219 
* OUTPUT: br_219 
* OUTPUT: bl_220 
* OUTPUT: br_220 
* OUTPUT: bl_221 
* OUTPUT: br_221 
* OUTPUT: bl_222 
* OUTPUT: br_222 
* OUTPUT: bl_223 
* OUTPUT: br_223 
* OUTPUT: bl_224 
* OUTPUT: br_224 
* OUTPUT: bl_225 
* OUTPUT: br_225 
* OUTPUT: bl_226 
* OUTPUT: br_226 
* OUTPUT: bl_227 
* OUTPUT: br_227 
* OUTPUT: bl_228 
* OUTPUT: br_228 
* OUTPUT: bl_229 
* OUTPUT: br_229 
* OUTPUT: bl_230 
* OUTPUT: br_230 
* OUTPUT: bl_231 
* OUTPUT: br_231 
* OUTPUT: bl_232 
* OUTPUT: br_232 
* OUTPUT: bl_233 
* OUTPUT: br_233 
* OUTPUT: bl_234 
* OUTPUT: br_234 
* OUTPUT: bl_235 
* OUTPUT: br_235 
* OUTPUT: bl_236 
* OUTPUT: br_236 
* OUTPUT: bl_237 
* OUTPUT: br_237 
* OUTPUT: bl_238 
* OUTPUT: br_238 
* OUTPUT: bl_239 
* OUTPUT: br_239 
* OUTPUT: bl_240 
* OUTPUT: br_240 
* OUTPUT: bl_241 
* OUTPUT: br_241 
* OUTPUT: bl_242 
* OUTPUT: br_242 
* OUTPUT: bl_243 
* OUTPUT: br_243 
* OUTPUT: bl_244 
* OUTPUT: br_244 
* OUTPUT: bl_245 
* OUTPUT: br_245 
* OUTPUT: bl_246 
* OUTPUT: br_246 
* OUTPUT: bl_247 
* OUTPUT: br_247 
* OUTPUT: bl_248 
* OUTPUT: br_248 
* OUTPUT: bl_249 
* OUTPUT: br_249 
* OUTPUT: bl_250 
* OUTPUT: br_250 
* OUTPUT: bl_251 
* OUTPUT: br_251 
* OUTPUT: bl_252 
* OUTPUT: br_252 
* OUTPUT: bl_253 
* OUTPUT: br_253 
* OUTPUT: bl_254 
* OUTPUT: br_254 
* OUTPUT: bl_255 
* OUTPUT: br_255 
* OUTPUT: bl_256 
* OUTPUT: br_256 
* INPUT : en_bar 
* POWER : vdd 
* cols: 257 size: 1 bl: bl br: br
Xpre_column_0
+ bl_0 br_0 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_1
+ bl_1 br_1 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_2
+ bl_2 br_2 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_3
+ bl_3 br_3 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_4
+ bl_4 br_4 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_5
+ bl_5 br_5 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_6
+ bl_6 br_6 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_7
+ bl_7 br_7 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_8
+ bl_8 br_8 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_9
+ bl_9 br_9 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_10
+ bl_10 br_10 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_11
+ bl_11 br_11 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_12
+ bl_12 br_12 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_13
+ bl_13 br_13 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_14
+ bl_14 br_14 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_15
+ bl_15 br_15 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_16
+ bl_16 br_16 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_17
+ bl_17 br_17 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_18
+ bl_18 br_18 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_19
+ bl_19 br_19 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_20
+ bl_20 br_20 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_21
+ bl_21 br_21 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_22
+ bl_22 br_22 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_23
+ bl_23 br_23 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_24
+ bl_24 br_24 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_25
+ bl_25 br_25 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_26
+ bl_26 br_26 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_27
+ bl_27 br_27 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_28
+ bl_28 br_28 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_29
+ bl_29 br_29 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_30
+ bl_30 br_30 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_31
+ bl_31 br_31 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_32
+ bl_32 br_32 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_33
+ bl_33 br_33 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_34
+ bl_34 br_34 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_35
+ bl_35 br_35 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_36
+ bl_36 br_36 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_37
+ bl_37 br_37 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_38
+ bl_38 br_38 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_39
+ bl_39 br_39 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_40
+ bl_40 br_40 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_41
+ bl_41 br_41 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_42
+ bl_42 br_42 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_43
+ bl_43 br_43 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_44
+ bl_44 br_44 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_45
+ bl_45 br_45 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_46
+ bl_46 br_46 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_47
+ bl_47 br_47 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_48
+ bl_48 br_48 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_49
+ bl_49 br_49 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_50
+ bl_50 br_50 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_51
+ bl_51 br_51 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_52
+ bl_52 br_52 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_53
+ bl_53 br_53 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_54
+ bl_54 br_54 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_55
+ bl_55 br_55 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_56
+ bl_56 br_56 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_57
+ bl_57 br_57 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_58
+ bl_58 br_58 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_59
+ bl_59 br_59 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_60
+ bl_60 br_60 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_61
+ bl_61 br_61 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_62
+ bl_62 br_62 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_63
+ bl_63 br_63 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_64
+ bl_64 br_64 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_65
+ bl_65 br_65 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_66
+ bl_66 br_66 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_67
+ bl_67 br_67 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_68
+ bl_68 br_68 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_69
+ bl_69 br_69 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_70
+ bl_70 br_70 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_71
+ bl_71 br_71 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_72
+ bl_72 br_72 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_73
+ bl_73 br_73 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_74
+ bl_74 br_74 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_75
+ bl_75 br_75 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_76
+ bl_76 br_76 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_77
+ bl_77 br_77 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_78
+ bl_78 br_78 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_79
+ bl_79 br_79 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_80
+ bl_80 br_80 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_81
+ bl_81 br_81 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_82
+ bl_82 br_82 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_83
+ bl_83 br_83 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_84
+ bl_84 br_84 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_85
+ bl_85 br_85 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_86
+ bl_86 br_86 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_87
+ bl_87 br_87 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_88
+ bl_88 br_88 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_89
+ bl_89 br_89 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_90
+ bl_90 br_90 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_91
+ bl_91 br_91 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_92
+ bl_92 br_92 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_93
+ bl_93 br_93 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_94
+ bl_94 br_94 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_95
+ bl_95 br_95 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_96
+ bl_96 br_96 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_97
+ bl_97 br_97 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_98
+ bl_98 br_98 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_99
+ bl_99 br_99 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_100
+ bl_100 br_100 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_101
+ bl_101 br_101 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_102
+ bl_102 br_102 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_103
+ bl_103 br_103 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_104
+ bl_104 br_104 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_105
+ bl_105 br_105 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_106
+ bl_106 br_106 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_107
+ bl_107 br_107 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_108
+ bl_108 br_108 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_109
+ bl_109 br_109 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_110
+ bl_110 br_110 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_111
+ bl_111 br_111 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_112
+ bl_112 br_112 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_113
+ bl_113 br_113 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_114
+ bl_114 br_114 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_115
+ bl_115 br_115 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_116
+ bl_116 br_116 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_117
+ bl_117 br_117 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_118
+ bl_118 br_118 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_119
+ bl_119 br_119 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_120
+ bl_120 br_120 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_121
+ bl_121 br_121 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_122
+ bl_122 br_122 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_123
+ bl_123 br_123 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_124
+ bl_124 br_124 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_125
+ bl_125 br_125 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_126
+ bl_126 br_126 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_127
+ bl_127 br_127 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_128
+ bl_128 br_128 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_129
+ bl_129 br_129 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_130
+ bl_130 br_130 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_131
+ bl_131 br_131 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_132
+ bl_132 br_132 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_133
+ bl_133 br_133 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_134
+ bl_134 br_134 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_135
+ bl_135 br_135 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_136
+ bl_136 br_136 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_137
+ bl_137 br_137 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_138
+ bl_138 br_138 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_139
+ bl_139 br_139 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_140
+ bl_140 br_140 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_141
+ bl_141 br_141 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_142
+ bl_142 br_142 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_143
+ bl_143 br_143 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_144
+ bl_144 br_144 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_145
+ bl_145 br_145 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_146
+ bl_146 br_146 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_147
+ bl_147 br_147 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_148
+ bl_148 br_148 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_149
+ bl_149 br_149 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_150
+ bl_150 br_150 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_151
+ bl_151 br_151 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_152
+ bl_152 br_152 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_153
+ bl_153 br_153 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_154
+ bl_154 br_154 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_155
+ bl_155 br_155 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_156
+ bl_156 br_156 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_157
+ bl_157 br_157 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_158
+ bl_158 br_158 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_159
+ bl_159 br_159 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_160
+ bl_160 br_160 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_161
+ bl_161 br_161 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_162
+ bl_162 br_162 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_163
+ bl_163 br_163 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_164
+ bl_164 br_164 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_165
+ bl_165 br_165 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_166
+ bl_166 br_166 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_167
+ bl_167 br_167 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_168
+ bl_168 br_168 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_169
+ bl_169 br_169 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_170
+ bl_170 br_170 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_171
+ bl_171 br_171 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_172
+ bl_172 br_172 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_173
+ bl_173 br_173 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_174
+ bl_174 br_174 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_175
+ bl_175 br_175 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_176
+ bl_176 br_176 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_177
+ bl_177 br_177 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_178
+ bl_178 br_178 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_179
+ bl_179 br_179 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_180
+ bl_180 br_180 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_181
+ bl_181 br_181 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_182
+ bl_182 br_182 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_183
+ bl_183 br_183 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_184
+ bl_184 br_184 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_185
+ bl_185 br_185 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_186
+ bl_186 br_186 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_187
+ bl_187 br_187 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_188
+ bl_188 br_188 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_189
+ bl_189 br_189 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_190
+ bl_190 br_190 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_191
+ bl_191 br_191 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_192
+ bl_192 br_192 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_193
+ bl_193 br_193 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_194
+ bl_194 br_194 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_195
+ bl_195 br_195 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_196
+ bl_196 br_196 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_197
+ bl_197 br_197 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_198
+ bl_198 br_198 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_199
+ bl_199 br_199 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_200
+ bl_200 br_200 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_201
+ bl_201 br_201 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_202
+ bl_202 br_202 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_203
+ bl_203 br_203 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_204
+ bl_204 br_204 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_205
+ bl_205 br_205 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_206
+ bl_206 br_206 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_207
+ bl_207 br_207 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_208
+ bl_208 br_208 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_209
+ bl_209 br_209 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_210
+ bl_210 br_210 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_211
+ bl_211 br_211 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_212
+ bl_212 br_212 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_213
+ bl_213 br_213 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_214
+ bl_214 br_214 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_215
+ bl_215 br_215 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_216
+ bl_216 br_216 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_217
+ bl_217 br_217 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_218
+ bl_218 br_218 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_219
+ bl_219 br_219 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_220
+ bl_220 br_220 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_221
+ bl_221 br_221 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_222
+ bl_222 br_222 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_223
+ bl_223 br_223 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_224
+ bl_224 br_224 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_225
+ bl_225 br_225 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_226
+ bl_226 br_226 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_227
+ bl_227 br_227 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_228
+ bl_228 br_228 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_229
+ bl_229 br_229 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_230
+ bl_230 br_230 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_231
+ bl_231 br_231 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_232
+ bl_232 br_232 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_233
+ bl_233 br_233 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_234
+ bl_234 br_234 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_235
+ bl_235 br_235 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_236
+ bl_236 br_236 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_237
+ bl_237 br_237 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_238
+ bl_238 br_238 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_239
+ bl_239 br_239 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_240
+ bl_240 br_240 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_241
+ bl_241 br_241 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_242
+ bl_242 br_242 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_243
+ bl_243 br_243 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_244
+ bl_244 br_244 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_245
+ bl_245 br_245 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_246
+ bl_246 br_246 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_247
+ bl_247 br_247 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_248
+ bl_248 br_248 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_249
+ bl_249 br_249 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_250
+ bl_250 br_250 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_251
+ bl_251 br_251 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_252
+ bl_252 br_252 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_253
+ bl_253 br_253 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_254
+ bl_254 br_254 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_255
+ bl_255 br_255 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
Xpre_column_256
+ bl_256 br_256 en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_0
.ENDS sram_1rw0r0w_32_1024_freepdk45_precharge_array

.SUBCKT sense_amp bl br dout en vdd gnd
M_1 dint net_1 vdd vdd pmos_vtg w=540.0n l=50.0n
M_3 net_1 dint vdd vdd pmos_vtg w=540.0n l=50.0n
M_2 dint net_1 net_2 gnd nmos_vtg w=270.0n l=50.0n
M_8 net_1 dint net_2 gnd nmos_vtg w=270.0n l=50.0n
M_5 bl en dint vdd pmos_vtg w=720.0n l=50.0n
M_6 br en net_1 vdd pmos_vtg w=720.0n l=50.0n
M_7 net_2 en gnd gnd nmos_vtg w=270.0n l=50.0n

M_9 dout_bar dint vdd vdd pmos_vtg w=180.0n l=50.0n
M_10 dout_bar dint gnd gnd nmos_vtg w=90.0n l=50.0n
M_11 dout dout_bar vdd vdd pmos_vtg w=540.0n l=50.0n
M_12 dout dout_bar gnd gnd nmos_vtg w=270.0n l=50.0n
.ENDS sense_amp


.SUBCKT sram_1rw0r0w_32_1024_freepdk45_sense_amp_array
+ data_0 bl_0 br_0 data_1 bl_1 br_1 data_2 bl_2 br_2 data_3 bl_3 br_3
+ data_4 bl_4 br_4 data_5 bl_5 br_5 data_6 bl_6 br_6 data_7 bl_7 br_7
+ data_8 bl_8 br_8 data_9 bl_9 br_9 data_10 bl_10 br_10 data_11 bl_11
+ br_11 data_12 bl_12 br_12 data_13 bl_13 br_13 data_14 bl_14 br_14
+ data_15 bl_15 br_15 data_16 bl_16 br_16 data_17 bl_17 br_17 data_18
+ bl_18 br_18 data_19 bl_19 br_19 data_20 bl_20 br_20 data_21 bl_21
+ br_21 data_22 bl_22 br_22 data_23 bl_23 br_23 data_24 bl_24 br_24
+ data_25 bl_25 br_25 data_26 bl_26 br_26 data_27 bl_27 br_27 data_28
+ bl_28 br_28 data_29 bl_29 br_29 data_30 bl_30 br_30 data_31 bl_31
+ br_31 en vdd gnd
* OUTPUT: data_0 
* INPUT : bl_0 
* INPUT : br_0 
* OUTPUT: data_1 
* INPUT : bl_1 
* INPUT : br_1 
* OUTPUT: data_2 
* INPUT : bl_2 
* INPUT : br_2 
* OUTPUT: data_3 
* INPUT : bl_3 
* INPUT : br_3 
* OUTPUT: data_4 
* INPUT : bl_4 
* INPUT : br_4 
* OUTPUT: data_5 
* INPUT : bl_5 
* INPUT : br_5 
* OUTPUT: data_6 
* INPUT : bl_6 
* INPUT : br_6 
* OUTPUT: data_7 
* INPUT : bl_7 
* INPUT : br_7 
* OUTPUT: data_8 
* INPUT : bl_8 
* INPUT : br_8 
* OUTPUT: data_9 
* INPUT : bl_9 
* INPUT : br_9 
* OUTPUT: data_10 
* INPUT : bl_10 
* INPUT : br_10 
* OUTPUT: data_11 
* INPUT : bl_11 
* INPUT : br_11 
* OUTPUT: data_12 
* INPUT : bl_12 
* INPUT : br_12 
* OUTPUT: data_13 
* INPUT : bl_13 
* INPUT : br_13 
* OUTPUT: data_14 
* INPUT : bl_14 
* INPUT : br_14 
* OUTPUT: data_15 
* INPUT : bl_15 
* INPUT : br_15 
* OUTPUT: data_16 
* INPUT : bl_16 
* INPUT : br_16 
* OUTPUT: data_17 
* INPUT : bl_17 
* INPUT : br_17 
* OUTPUT: data_18 
* INPUT : bl_18 
* INPUT : br_18 
* OUTPUT: data_19 
* INPUT : bl_19 
* INPUT : br_19 
* OUTPUT: data_20 
* INPUT : bl_20 
* INPUT : br_20 
* OUTPUT: data_21 
* INPUT : bl_21 
* INPUT : br_21 
* OUTPUT: data_22 
* INPUT : bl_22 
* INPUT : br_22 
* OUTPUT: data_23 
* INPUT : bl_23 
* INPUT : br_23 
* OUTPUT: data_24 
* INPUT : bl_24 
* INPUT : br_24 
* OUTPUT: data_25 
* INPUT : bl_25 
* INPUT : br_25 
* OUTPUT: data_26 
* INPUT : bl_26 
* INPUT : br_26 
* OUTPUT: data_27 
* INPUT : bl_27 
* INPUT : br_27 
* OUTPUT: data_28 
* INPUT : bl_28 
* INPUT : br_28 
* OUTPUT: data_29 
* INPUT : bl_29 
* INPUT : br_29 
* OUTPUT: data_30 
* INPUT : bl_30 
* INPUT : br_30 
* OUTPUT: data_31 
* INPUT : bl_31 
* INPUT : br_31 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* word_size 32
* words_per_row: 8
Xsa_d0
+ bl_0 br_0 data_0 en vdd gnd
+ sense_amp
Xsa_d1
+ bl_1 br_1 data_1 en vdd gnd
+ sense_amp
Xsa_d2
+ bl_2 br_2 data_2 en vdd gnd
+ sense_amp
Xsa_d3
+ bl_3 br_3 data_3 en vdd gnd
+ sense_amp
Xsa_d4
+ bl_4 br_4 data_4 en vdd gnd
+ sense_amp
Xsa_d5
+ bl_5 br_5 data_5 en vdd gnd
+ sense_amp
Xsa_d6
+ bl_6 br_6 data_6 en vdd gnd
+ sense_amp
Xsa_d7
+ bl_7 br_7 data_7 en vdd gnd
+ sense_amp
Xsa_d8
+ bl_8 br_8 data_8 en vdd gnd
+ sense_amp
Xsa_d9
+ bl_9 br_9 data_9 en vdd gnd
+ sense_amp
Xsa_d10
+ bl_10 br_10 data_10 en vdd gnd
+ sense_amp
Xsa_d11
+ bl_11 br_11 data_11 en vdd gnd
+ sense_amp
Xsa_d12
+ bl_12 br_12 data_12 en vdd gnd
+ sense_amp
Xsa_d13
+ bl_13 br_13 data_13 en vdd gnd
+ sense_amp
Xsa_d14
+ bl_14 br_14 data_14 en vdd gnd
+ sense_amp
Xsa_d15
+ bl_15 br_15 data_15 en vdd gnd
+ sense_amp
Xsa_d16
+ bl_16 br_16 data_16 en vdd gnd
+ sense_amp
Xsa_d17
+ bl_17 br_17 data_17 en vdd gnd
+ sense_amp
Xsa_d18
+ bl_18 br_18 data_18 en vdd gnd
+ sense_amp
Xsa_d19
+ bl_19 br_19 data_19 en vdd gnd
+ sense_amp
Xsa_d20
+ bl_20 br_20 data_20 en vdd gnd
+ sense_amp
Xsa_d21
+ bl_21 br_21 data_21 en vdd gnd
+ sense_amp
Xsa_d22
+ bl_22 br_22 data_22 en vdd gnd
+ sense_amp
Xsa_d23
+ bl_23 br_23 data_23 en vdd gnd
+ sense_amp
Xsa_d24
+ bl_24 br_24 data_24 en vdd gnd
+ sense_amp
Xsa_d25
+ bl_25 br_25 data_25 en vdd gnd
+ sense_amp
Xsa_d26
+ bl_26 br_26 data_26 en vdd gnd
+ sense_amp
Xsa_d27
+ bl_27 br_27 data_27 en vdd gnd
+ sense_amp
Xsa_d28
+ bl_28 br_28 data_28 en vdd gnd
+ sense_amp
Xsa_d29
+ bl_29 br_29 data_29 en vdd gnd
+ sense_amp
Xsa_d30
+ bl_30 br_30 data_30 en vdd gnd
+ sense_amp
Xsa_d31
+ bl_31 br_31 data_31 en vdd gnd
+ sense_amp
.ENDS sram_1rw0r0w_32_1024_freepdk45_sense_amp_array

* spice ptx M{0} {1} nmos_vtg m=1 w=0.72u l=0.05u pd=1.54u ps=1.54u as=0.09p ad=0.09p

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_column_mux
+ bl br bl_out br_out sel gnd
* INOUT : bl 
* INOUT : br 
* INOUT : bl_out 
* INOUT : br_out 
* INOUT : sel 
* INOUT : gnd 
Mmux_tx1 bl sel bl_out gnd nmos_vtg m=1 w=0.72u l=0.05u pd=1.54u ps=1.54u as=0.09p ad=0.09p
Mmux_tx2 br sel br_out gnd nmos_vtg m=1 w=0.72u l=0.05u pd=1.54u ps=1.54u as=0.09p ad=0.09p
.ENDS sram_1rw0r0w_32_1024_freepdk45_column_mux

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_column_mux_array
+ bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6
+ bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12
+ bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18
+ br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23
+ bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29
+ br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34
+ bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40
+ br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45
+ bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51
+ br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56
+ bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62
+ br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67
+ bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73
+ br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78
+ bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84
+ br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89
+ bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95
+ br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100
+ bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105
+ bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110
+ bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115
+ bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120
+ bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125
+ bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130
+ bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135
+ bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140
+ bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145
+ bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150
+ bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155
+ bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160
+ bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165
+ bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170
+ bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175
+ bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180
+ bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185
+ bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190
+ bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195
+ bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200
+ bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205
+ bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210
+ bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215
+ bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220
+ bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225
+ bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230
+ bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235
+ bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240
+ bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245
+ bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250
+ bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255
+ sel_0 sel_1 sel_2 sel_3 sel_4 sel_5 sel_6 sel_7 bl_out_0 br_out_0
+ bl_out_1 br_out_1 bl_out_2 br_out_2 bl_out_3 br_out_3 bl_out_4
+ br_out_4 bl_out_5 br_out_5 bl_out_6 br_out_6 bl_out_7 br_out_7
+ bl_out_8 br_out_8 bl_out_9 br_out_9 bl_out_10 br_out_10 bl_out_11
+ br_out_11 bl_out_12 br_out_12 bl_out_13 br_out_13 bl_out_14 br_out_14
+ bl_out_15 br_out_15 bl_out_16 br_out_16 bl_out_17 br_out_17 bl_out_18
+ br_out_18 bl_out_19 br_out_19 bl_out_20 br_out_20 bl_out_21 br_out_21
+ bl_out_22 br_out_22 bl_out_23 br_out_23 bl_out_24 br_out_24 bl_out_25
+ br_out_25 bl_out_26 br_out_26 bl_out_27 br_out_27 bl_out_28 br_out_28
+ bl_out_29 br_out_29 bl_out_30 br_out_30 bl_out_31 br_out_31 gnd
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : bl_64 
* INOUT : br_64 
* INOUT : bl_65 
* INOUT : br_65 
* INOUT : bl_66 
* INOUT : br_66 
* INOUT : bl_67 
* INOUT : br_67 
* INOUT : bl_68 
* INOUT : br_68 
* INOUT : bl_69 
* INOUT : br_69 
* INOUT : bl_70 
* INOUT : br_70 
* INOUT : bl_71 
* INOUT : br_71 
* INOUT : bl_72 
* INOUT : br_72 
* INOUT : bl_73 
* INOUT : br_73 
* INOUT : bl_74 
* INOUT : br_74 
* INOUT : bl_75 
* INOUT : br_75 
* INOUT : bl_76 
* INOUT : br_76 
* INOUT : bl_77 
* INOUT : br_77 
* INOUT : bl_78 
* INOUT : br_78 
* INOUT : bl_79 
* INOUT : br_79 
* INOUT : bl_80 
* INOUT : br_80 
* INOUT : bl_81 
* INOUT : br_81 
* INOUT : bl_82 
* INOUT : br_82 
* INOUT : bl_83 
* INOUT : br_83 
* INOUT : bl_84 
* INOUT : br_84 
* INOUT : bl_85 
* INOUT : br_85 
* INOUT : bl_86 
* INOUT : br_86 
* INOUT : bl_87 
* INOUT : br_87 
* INOUT : bl_88 
* INOUT : br_88 
* INOUT : bl_89 
* INOUT : br_89 
* INOUT : bl_90 
* INOUT : br_90 
* INOUT : bl_91 
* INOUT : br_91 
* INOUT : bl_92 
* INOUT : br_92 
* INOUT : bl_93 
* INOUT : br_93 
* INOUT : bl_94 
* INOUT : br_94 
* INOUT : bl_95 
* INOUT : br_95 
* INOUT : bl_96 
* INOUT : br_96 
* INOUT : bl_97 
* INOUT : br_97 
* INOUT : bl_98 
* INOUT : br_98 
* INOUT : bl_99 
* INOUT : br_99 
* INOUT : bl_100 
* INOUT : br_100 
* INOUT : bl_101 
* INOUT : br_101 
* INOUT : bl_102 
* INOUT : br_102 
* INOUT : bl_103 
* INOUT : br_103 
* INOUT : bl_104 
* INOUT : br_104 
* INOUT : bl_105 
* INOUT : br_105 
* INOUT : bl_106 
* INOUT : br_106 
* INOUT : bl_107 
* INOUT : br_107 
* INOUT : bl_108 
* INOUT : br_108 
* INOUT : bl_109 
* INOUT : br_109 
* INOUT : bl_110 
* INOUT : br_110 
* INOUT : bl_111 
* INOUT : br_111 
* INOUT : bl_112 
* INOUT : br_112 
* INOUT : bl_113 
* INOUT : br_113 
* INOUT : bl_114 
* INOUT : br_114 
* INOUT : bl_115 
* INOUT : br_115 
* INOUT : bl_116 
* INOUT : br_116 
* INOUT : bl_117 
* INOUT : br_117 
* INOUT : bl_118 
* INOUT : br_118 
* INOUT : bl_119 
* INOUT : br_119 
* INOUT : bl_120 
* INOUT : br_120 
* INOUT : bl_121 
* INOUT : br_121 
* INOUT : bl_122 
* INOUT : br_122 
* INOUT : bl_123 
* INOUT : br_123 
* INOUT : bl_124 
* INOUT : br_124 
* INOUT : bl_125 
* INOUT : br_125 
* INOUT : bl_126 
* INOUT : br_126 
* INOUT : bl_127 
* INOUT : br_127 
* INOUT : bl_128 
* INOUT : br_128 
* INOUT : bl_129 
* INOUT : br_129 
* INOUT : bl_130 
* INOUT : br_130 
* INOUT : bl_131 
* INOUT : br_131 
* INOUT : bl_132 
* INOUT : br_132 
* INOUT : bl_133 
* INOUT : br_133 
* INOUT : bl_134 
* INOUT : br_134 
* INOUT : bl_135 
* INOUT : br_135 
* INOUT : bl_136 
* INOUT : br_136 
* INOUT : bl_137 
* INOUT : br_137 
* INOUT : bl_138 
* INOUT : br_138 
* INOUT : bl_139 
* INOUT : br_139 
* INOUT : bl_140 
* INOUT : br_140 
* INOUT : bl_141 
* INOUT : br_141 
* INOUT : bl_142 
* INOUT : br_142 
* INOUT : bl_143 
* INOUT : br_143 
* INOUT : bl_144 
* INOUT : br_144 
* INOUT : bl_145 
* INOUT : br_145 
* INOUT : bl_146 
* INOUT : br_146 
* INOUT : bl_147 
* INOUT : br_147 
* INOUT : bl_148 
* INOUT : br_148 
* INOUT : bl_149 
* INOUT : br_149 
* INOUT : bl_150 
* INOUT : br_150 
* INOUT : bl_151 
* INOUT : br_151 
* INOUT : bl_152 
* INOUT : br_152 
* INOUT : bl_153 
* INOUT : br_153 
* INOUT : bl_154 
* INOUT : br_154 
* INOUT : bl_155 
* INOUT : br_155 
* INOUT : bl_156 
* INOUT : br_156 
* INOUT : bl_157 
* INOUT : br_157 
* INOUT : bl_158 
* INOUT : br_158 
* INOUT : bl_159 
* INOUT : br_159 
* INOUT : bl_160 
* INOUT : br_160 
* INOUT : bl_161 
* INOUT : br_161 
* INOUT : bl_162 
* INOUT : br_162 
* INOUT : bl_163 
* INOUT : br_163 
* INOUT : bl_164 
* INOUT : br_164 
* INOUT : bl_165 
* INOUT : br_165 
* INOUT : bl_166 
* INOUT : br_166 
* INOUT : bl_167 
* INOUT : br_167 
* INOUT : bl_168 
* INOUT : br_168 
* INOUT : bl_169 
* INOUT : br_169 
* INOUT : bl_170 
* INOUT : br_170 
* INOUT : bl_171 
* INOUT : br_171 
* INOUT : bl_172 
* INOUT : br_172 
* INOUT : bl_173 
* INOUT : br_173 
* INOUT : bl_174 
* INOUT : br_174 
* INOUT : bl_175 
* INOUT : br_175 
* INOUT : bl_176 
* INOUT : br_176 
* INOUT : bl_177 
* INOUT : br_177 
* INOUT : bl_178 
* INOUT : br_178 
* INOUT : bl_179 
* INOUT : br_179 
* INOUT : bl_180 
* INOUT : br_180 
* INOUT : bl_181 
* INOUT : br_181 
* INOUT : bl_182 
* INOUT : br_182 
* INOUT : bl_183 
* INOUT : br_183 
* INOUT : bl_184 
* INOUT : br_184 
* INOUT : bl_185 
* INOUT : br_185 
* INOUT : bl_186 
* INOUT : br_186 
* INOUT : bl_187 
* INOUT : br_187 
* INOUT : bl_188 
* INOUT : br_188 
* INOUT : bl_189 
* INOUT : br_189 
* INOUT : bl_190 
* INOUT : br_190 
* INOUT : bl_191 
* INOUT : br_191 
* INOUT : bl_192 
* INOUT : br_192 
* INOUT : bl_193 
* INOUT : br_193 
* INOUT : bl_194 
* INOUT : br_194 
* INOUT : bl_195 
* INOUT : br_195 
* INOUT : bl_196 
* INOUT : br_196 
* INOUT : bl_197 
* INOUT : br_197 
* INOUT : bl_198 
* INOUT : br_198 
* INOUT : bl_199 
* INOUT : br_199 
* INOUT : bl_200 
* INOUT : br_200 
* INOUT : bl_201 
* INOUT : br_201 
* INOUT : bl_202 
* INOUT : br_202 
* INOUT : bl_203 
* INOUT : br_203 
* INOUT : bl_204 
* INOUT : br_204 
* INOUT : bl_205 
* INOUT : br_205 
* INOUT : bl_206 
* INOUT : br_206 
* INOUT : bl_207 
* INOUT : br_207 
* INOUT : bl_208 
* INOUT : br_208 
* INOUT : bl_209 
* INOUT : br_209 
* INOUT : bl_210 
* INOUT : br_210 
* INOUT : bl_211 
* INOUT : br_211 
* INOUT : bl_212 
* INOUT : br_212 
* INOUT : bl_213 
* INOUT : br_213 
* INOUT : bl_214 
* INOUT : br_214 
* INOUT : bl_215 
* INOUT : br_215 
* INOUT : bl_216 
* INOUT : br_216 
* INOUT : bl_217 
* INOUT : br_217 
* INOUT : bl_218 
* INOUT : br_218 
* INOUT : bl_219 
* INOUT : br_219 
* INOUT : bl_220 
* INOUT : br_220 
* INOUT : bl_221 
* INOUT : br_221 
* INOUT : bl_222 
* INOUT : br_222 
* INOUT : bl_223 
* INOUT : br_223 
* INOUT : bl_224 
* INOUT : br_224 
* INOUT : bl_225 
* INOUT : br_225 
* INOUT : bl_226 
* INOUT : br_226 
* INOUT : bl_227 
* INOUT : br_227 
* INOUT : bl_228 
* INOUT : br_228 
* INOUT : bl_229 
* INOUT : br_229 
* INOUT : bl_230 
* INOUT : br_230 
* INOUT : bl_231 
* INOUT : br_231 
* INOUT : bl_232 
* INOUT : br_232 
* INOUT : bl_233 
* INOUT : br_233 
* INOUT : bl_234 
* INOUT : br_234 
* INOUT : bl_235 
* INOUT : br_235 
* INOUT : bl_236 
* INOUT : br_236 
* INOUT : bl_237 
* INOUT : br_237 
* INOUT : bl_238 
* INOUT : br_238 
* INOUT : bl_239 
* INOUT : br_239 
* INOUT : bl_240 
* INOUT : br_240 
* INOUT : bl_241 
* INOUT : br_241 
* INOUT : bl_242 
* INOUT : br_242 
* INOUT : bl_243 
* INOUT : br_243 
* INOUT : bl_244 
* INOUT : br_244 
* INOUT : bl_245 
* INOUT : br_245 
* INOUT : bl_246 
* INOUT : br_246 
* INOUT : bl_247 
* INOUT : br_247 
* INOUT : bl_248 
* INOUT : br_248 
* INOUT : bl_249 
* INOUT : br_249 
* INOUT : bl_250 
* INOUT : br_250 
* INOUT : bl_251 
* INOUT : br_251 
* INOUT : bl_252 
* INOUT : br_252 
* INOUT : bl_253 
* INOUT : br_253 
* INOUT : bl_254 
* INOUT : br_254 
* INOUT : bl_255 
* INOUT : br_255 
* INOUT : sel_0 
* INOUT : sel_1 
* INOUT : sel_2 
* INOUT : sel_3 
* INOUT : sel_4 
* INOUT : sel_5 
* INOUT : sel_6 
* INOUT : sel_7 
* INOUT : bl_out_0 
* INOUT : br_out_0 
* INOUT : bl_out_1 
* INOUT : br_out_1 
* INOUT : bl_out_2 
* INOUT : br_out_2 
* INOUT : bl_out_3 
* INOUT : br_out_3 
* INOUT : bl_out_4 
* INOUT : br_out_4 
* INOUT : bl_out_5 
* INOUT : br_out_5 
* INOUT : bl_out_6 
* INOUT : br_out_6 
* INOUT : bl_out_7 
* INOUT : br_out_7 
* INOUT : bl_out_8 
* INOUT : br_out_8 
* INOUT : bl_out_9 
* INOUT : br_out_9 
* INOUT : bl_out_10 
* INOUT : br_out_10 
* INOUT : bl_out_11 
* INOUT : br_out_11 
* INOUT : bl_out_12 
* INOUT : br_out_12 
* INOUT : bl_out_13 
* INOUT : br_out_13 
* INOUT : bl_out_14 
* INOUT : br_out_14 
* INOUT : bl_out_15 
* INOUT : br_out_15 
* INOUT : bl_out_16 
* INOUT : br_out_16 
* INOUT : bl_out_17 
* INOUT : br_out_17 
* INOUT : bl_out_18 
* INOUT : br_out_18 
* INOUT : bl_out_19 
* INOUT : br_out_19 
* INOUT : bl_out_20 
* INOUT : br_out_20 
* INOUT : bl_out_21 
* INOUT : br_out_21 
* INOUT : bl_out_22 
* INOUT : br_out_22 
* INOUT : bl_out_23 
* INOUT : br_out_23 
* INOUT : bl_out_24 
* INOUT : br_out_24 
* INOUT : bl_out_25 
* INOUT : br_out_25 
* INOUT : bl_out_26 
* INOUT : br_out_26 
* INOUT : bl_out_27 
* INOUT : br_out_27 
* INOUT : bl_out_28 
* INOUT : br_out_28 
* INOUT : bl_out_29 
* INOUT : br_out_29 
* INOUT : bl_out_30 
* INOUT : br_out_30 
* INOUT : bl_out_31 
* INOUT : br_out_31 
* INOUT : gnd 
* cols: 256 word_size: 32 bl: bl br: br
XXMUX0
+ bl_0 br_0 bl_out_0 br_out_0 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX1
+ bl_1 br_1 bl_out_0 br_out_0 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX2
+ bl_2 br_2 bl_out_0 br_out_0 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX3
+ bl_3 br_3 bl_out_0 br_out_0 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX4
+ bl_4 br_4 bl_out_0 br_out_0 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX5
+ bl_5 br_5 bl_out_0 br_out_0 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX6
+ bl_6 br_6 bl_out_0 br_out_0 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX7
+ bl_7 br_7 bl_out_0 br_out_0 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX8
+ bl_8 br_8 bl_out_1 br_out_1 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX9
+ bl_9 br_9 bl_out_1 br_out_1 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX10
+ bl_10 br_10 bl_out_1 br_out_1 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX11
+ bl_11 br_11 bl_out_1 br_out_1 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX12
+ bl_12 br_12 bl_out_1 br_out_1 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX13
+ bl_13 br_13 bl_out_1 br_out_1 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX14
+ bl_14 br_14 bl_out_1 br_out_1 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX15
+ bl_15 br_15 bl_out_1 br_out_1 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX16
+ bl_16 br_16 bl_out_2 br_out_2 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX17
+ bl_17 br_17 bl_out_2 br_out_2 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX18
+ bl_18 br_18 bl_out_2 br_out_2 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX19
+ bl_19 br_19 bl_out_2 br_out_2 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX20
+ bl_20 br_20 bl_out_2 br_out_2 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX21
+ bl_21 br_21 bl_out_2 br_out_2 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX22
+ bl_22 br_22 bl_out_2 br_out_2 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX23
+ bl_23 br_23 bl_out_2 br_out_2 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX24
+ bl_24 br_24 bl_out_3 br_out_3 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX25
+ bl_25 br_25 bl_out_3 br_out_3 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX26
+ bl_26 br_26 bl_out_3 br_out_3 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX27
+ bl_27 br_27 bl_out_3 br_out_3 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX28
+ bl_28 br_28 bl_out_3 br_out_3 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX29
+ bl_29 br_29 bl_out_3 br_out_3 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX30
+ bl_30 br_30 bl_out_3 br_out_3 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX31
+ bl_31 br_31 bl_out_3 br_out_3 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX32
+ bl_32 br_32 bl_out_4 br_out_4 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX33
+ bl_33 br_33 bl_out_4 br_out_4 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX34
+ bl_34 br_34 bl_out_4 br_out_4 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX35
+ bl_35 br_35 bl_out_4 br_out_4 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX36
+ bl_36 br_36 bl_out_4 br_out_4 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX37
+ bl_37 br_37 bl_out_4 br_out_4 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX38
+ bl_38 br_38 bl_out_4 br_out_4 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX39
+ bl_39 br_39 bl_out_4 br_out_4 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX40
+ bl_40 br_40 bl_out_5 br_out_5 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX41
+ bl_41 br_41 bl_out_5 br_out_5 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX42
+ bl_42 br_42 bl_out_5 br_out_5 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX43
+ bl_43 br_43 bl_out_5 br_out_5 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX44
+ bl_44 br_44 bl_out_5 br_out_5 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX45
+ bl_45 br_45 bl_out_5 br_out_5 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX46
+ bl_46 br_46 bl_out_5 br_out_5 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX47
+ bl_47 br_47 bl_out_5 br_out_5 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX48
+ bl_48 br_48 bl_out_6 br_out_6 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX49
+ bl_49 br_49 bl_out_6 br_out_6 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX50
+ bl_50 br_50 bl_out_6 br_out_6 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX51
+ bl_51 br_51 bl_out_6 br_out_6 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX52
+ bl_52 br_52 bl_out_6 br_out_6 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX53
+ bl_53 br_53 bl_out_6 br_out_6 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX54
+ bl_54 br_54 bl_out_6 br_out_6 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX55
+ bl_55 br_55 bl_out_6 br_out_6 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX56
+ bl_56 br_56 bl_out_7 br_out_7 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX57
+ bl_57 br_57 bl_out_7 br_out_7 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX58
+ bl_58 br_58 bl_out_7 br_out_7 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX59
+ bl_59 br_59 bl_out_7 br_out_7 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX60
+ bl_60 br_60 bl_out_7 br_out_7 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX61
+ bl_61 br_61 bl_out_7 br_out_7 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX62
+ bl_62 br_62 bl_out_7 br_out_7 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX63
+ bl_63 br_63 bl_out_7 br_out_7 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX64
+ bl_64 br_64 bl_out_8 br_out_8 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX65
+ bl_65 br_65 bl_out_8 br_out_8 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX66
+ bl_66 br_66 bl_out_8 br_out_8 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX67
+ bl_67 br_67 bl_out_8 br_out_8 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX68
+ bl_68 br_68 bl_out_8 br_out_8 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX69
+ bl_69 br_69 bl_out_8 br_out_8 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX70
+ bl_70 br_70 bl_out_8 br_out_8 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX71
+ bl_71 br_71 bl_out_8 br_out_8 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX72
+ bl_72 br_72 bl_out_9 br_out_9 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX73
+ bl_73 br_73 bl_out_9 br_out_9 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX74
+ bl_74 br_74 bl_out_9 br_out_9 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX75
+ bl_75 br_75 bl_out_9 br_out_9 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX76
+ bl_76 br_76 bl_out_9 br_out_9 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX77
+ bl_77 br_77 bl_out_9 br_out_9 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX78
+ bl_78 br_78 bl_out_9 br_out_9 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX79
+ bl_79 br_79 bl_out_9 br_out_9 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX80
+ bl_80 br_80 bl_out_10 br_out_10 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX81
+ bl_81 br_81 bl_out_10 br_out_10 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX82
+ bl_82 br_82 bl_out_10 br_out_10 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX83
+ bl_83 br_83 bl_out_10 br_out_10 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX84
+ bl_84 br_84 bl_out_10 br_out_10 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX85
+ bl_85 br_85 bl_out_10 br_out_10 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX86
+ bl_86 br_86 bl_out_10 br_out_10 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX87
+ bl_87 br_87 bl_out_10 br_out_10 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX88
+ bl_88 br_88 bl_out_11 br_out_11 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX89
+ bl_89 br_89 bl_out_11 br_out_11 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX90
+ bl_90 br_90 bl_out_11 br_out_11 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX91
+ bl_91 br_91 bl_out_11 br_out_11 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX92
+ bl_92 br_92 bl_out_11 br_out_11 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX93
+ bl_93 br_93 bl_out_11 br_out_11 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX94
+ bl_94 br_94 bl_out_11 br_out_11 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX95
+ bl_95 br_95 bl_out_11 br_out_11 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX96
+ bl_96 br_96 bl_out_12 br_out_12 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX97
+ bl_97 br_97 bl_out_12 br_out_12 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX98
+ bl_98 br_98 bl_out_12 br_out_12 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX99
+ bl_99 br_99 bl_out_12 br_out_12 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX100
+ bl_100 br_100 bl_out_12 br_out_12 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX101
+ bl_101 br_101 bl_out_12 br_out_12 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX102
+ bl_102 br_102 bl_out_12 br_out_12 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX103
+ bl_103 br_103 bl_out_12 br_out_12 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX104
+ bl_104 br_104 bl_out_13 br_out_13 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX105
+ bl_105 br_105 bl_out_13 br_out_13 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX106
+ bl_106 br_106 bl_out_13 br_out_13 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX107
+ bl_107 br_107 bl_out_13 br_out_13 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX108
+ bl_108 br_108 bl_out_13 br_out_13 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX109
+ bl_109 br_109 bl_out_13 br_out_13 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX110
+ bl_110 br_110 bl_out_13 br_out_13 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX111
+ bl_111 br_111 bl_out_13 br_out_13 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX112
+ bl_112 br_112 bl_out_14 br_out_14 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX113
+ bl_113 br_113 bl_out_14 br_out_14 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX114
+ bl_114 br_114 bl_out_14 br_out_14 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX115
+ bl_115 br_115 bl_out_14 br_out_14 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX116
+ bl_116 br_116 bl_out_14 br_out_14 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX117
+ bl_117 br_117 bl_out_14 br_out_14 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX118
+ bl_118 br_118 bl_out_14 br_out_14 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX119
+ bl_119 br_119 bl_out_14 br_out_14 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX120
+ bl_120 br_120 bl_out_15 br_out_15 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX121
+ bl_121 br_121 bl_out_15 br_out_15 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX122
+ bl_122 br_122 bl_out_15 br_out_15 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX123
+ bl_123 br_123 bl_out_15 br_out_15 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX124
+ bl_124 br_124 bl_out_15 br_out_15 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX125
+ bl_125 br_125 bl_out_15 br_out_15 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX126
+ bl_126 br_126 bl_out_15 br_out_15 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX127
+ bl_127 br_127 bl_out_15 br_out_15 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX128
+ bl_128 br_128 bl_out_16 br_out_16 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX129
+ bl_129 br_129 bl_out_16 br_out_16 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX130
+ bl_130 br_130 bl_out_16 br_out_16 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX131
+ bl_131 br_131 bl_out_16 br_out_16 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX132
+ bl_132 br_132 bl_out_16 br_out_16 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX133
+ bl_133 br_133 bl_out_16 br_out_16 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX134
+ bl_134 br_134 bl_out_16 br_out_16 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX135
+ bl_135 br_135 bl_out_16 br_out_16 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX136
+ bl_136 br_136 bl_out_17 br_out_17 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX137
+ bl_137 br_137 bl_out_17 br_out_17 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX138
+ bl_138 br_138 bl_out_17 br_out_17 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX139
+ bl_139 br_139 bl_out_17 br_out_17 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX140
+ bl_140 br_140 bl_out_17 br_out_17 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX141
+ bl_141 br_141 bl_out_17 br_out_17 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX142
+ bl_142 br_142 bl_out_17 br_out_17 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX143
+ bl_143 br_143 bl_out_17 br_out_17 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX144
+ bl_144 br_144 bl_out_18 br_out_18 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX145
+ bl_145 br_145 bl_out_18 br_out_18 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX146
+ bl_146 br_146 bl_out_18 br_out_18 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX147
+ bl_147 br_147 bl_out_18 br_out_18 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX148
+ bl_148 br_148 bl_out_18 br_out_18 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX149
+ bl_149 br_149 bl_out_18 br_out_18 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX150
+ bl_150 br_150 bl_out_18 br_out_18 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX151
+ bl_151 br_151 bl_out_18 br_out_18 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX152
+ bl_152 br_152 bl_out_19 br_out_19 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX153
+ bl_153 br_153 bl_out_19 br_out_19 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX154
+ bl_154 br_154 bl_out_19 br_out_19 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX155
+ bl_155 br_155 bl_out_19 br_out_19 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX156
+ bl_156 br_156 bl_out_19 br_out_19 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX157
+ bl_157 br_157 bl_out_19 br_out_19 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX158
+ bl_158 br_158 bl_out_19 br_out_19 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX159
+ bl_159 br_159 bl_out_19 br_out_19 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX160
+ bl_160 br_160 bl_out_20 br_out_20 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX161
+ bl_161 br_161 bl_out_20 br_out_20 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX162
+ bl_162 br_162 bl_out_20 br_out_20 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX163
+ bl_163 br_163 bl_out_20 br_out_20 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX164
+ bl_164 br_164 bl_out_20 br_out_20 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX165
+ bl_165 br_165 bl_out_20 br_out_20 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX166
+ bl_166 br_166 bl_out_20 br_out_20 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX167
+ bl_167 br_167 bl_out_20 br_out_20 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX168
+ bl_168 br_168 bl_out_21 br_out_21 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX169
+ bl_169 br_169 bl_out_21 br_out_21 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX170
+ bl_170 br_170 bl_out_21 br_out_21 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX171
+ bl_171 br_171 bl_out_21 br_out_21 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX172
+ bl_172 br_172 bl_out_21 br_out_21 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX173
+ bl_173 br_173 bl_out_21 br_out_21 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX174
+ bl_174 br_174 bl_out_21 br_out_21 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX175
+ bl_175 br_175 bl_out_21 br_out_21 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX176
+ bl_176 br_176 bl_out_22 br_out_22 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX177
+ bl_177 br_177 bl_out_22 br_out_22 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX178
+ bl_178 br_178 bl_out_22 br_out_22 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX179
+ bl_179 br_179 bl_out_22 br_out_22 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX180
+ bl_180 br_180 bl_out_22 br_out_22 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX181
+ bl_181 br_181 bl_out_22 br_out_22 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX182
+ bl_182 br_182 bl_out_22 br_out_22 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX183
+ bl_183 br_183 bl_out_22 br_out_22 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX184
+ bl_184 br_184 bl_out_23 br_out_23 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX185
+ bl_185 br_185 bl_out_23 br_out_23 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX186
+ bl_186 br_186 bl_out_23 br_out_23 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX187
+ bl_187 br_187 bl_out_23 br_out_23 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX188
+ bl_188 br_188 bl_out_23 br_out_23 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX189
+ bl_189 br_189 bl_out_23 br_out_23 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX190
+ bl_190 br_190 bl_out_23 br_out_23 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX191
+ bl_191 br_191 bl_out_23 br_out_23 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX192
+ bl_192 br_192 bl_out_24 br_out_24 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX193
+ bl_193 br_193 bl_out_24 br_out_24 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX194
+ bl_194 br_194 bl_out_24 br_out_24 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX195
+ bl_195 br_195 bl_out_24 br_out_24 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX196
+ bl_196 br_196 bl_out_24 br_out_24 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX197
+ bl_197 br_197 bl_out_24 br_out_24 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX198
+ bl_198 br_198 bl_out_24 br_out_24 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX199
+ bl_199 br_199 bl_out_24 br_out_24 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX200
+ bl_200 br_200 bl_out_25 br_out_25 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX201
+ bl_201 br_201 bl_out_25 br_out_25 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX202
+ bl_202 br_202 bl_out_25 br_out_25 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX203
+ bl_203 br_203 bl_out_25 br_out_25 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX204
+ bl_204 br_204 bl_out_25 br_out_25 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX205
+ bl_205 br_205 bl_out_25 br_out_25 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX206
+ bl_206 br_206 bl_out_25 br_out_25 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX207
+ bl_207 br_207 bl_out_25 br_out_25 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX208
+ bl_208 br_208 bl_out_26 br_out_26 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX209
+ bl_209 br_209 bl_out_26 br_out_26 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX210
+ bl_210 br_210 bl_out_26 br_out_26 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX211
+ bl_211 br_211 bl_out_26 br_out_26 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX212
+ bl_212 br_212 bl_out_26 br_out_26 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX213
+ bl_213 br_213 bl_out_26 br_out_26 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX214
+ bl_214 br_214 bl_out_26 br_out_26 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX215
+ bl_215 br_215 bl_out_26 br_out_26 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX216
+ bl_216 br_216 bl_out_27 br_out_27 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX217
+ bl_217 br_217 bl_out_27 br_out_27 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX218
+ bl_218 br_218 bl_out_27 br_out_27 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX219
+ bl_219 br_219 bl_out_27 br_out_27 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX220
+ bl_220 br_220 bl_out_27 br_out_27 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX221
+ bl_221 br_221 bl_out_27 br_out_27 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX222
+ bl_222 br_222 bl_out_27 br_out_27 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX223
+ bl_223 br_223 bl_out_27 br_out_27 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX224
+ bl_224 br_224 bl_out_28 br_out_28 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX225
+ bl_225 br_225 bl_out_28 br_out_28 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX226
+ bl_226 br_226 bl_out_28 br_out_28 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX227
+ bl_227 br_227 bl_out_28 br_out_28 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX228
+ bl_228 br_228 bl_out_28 br_out_28 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX229
+ bl_229 br_229 bl_out_28 br_out_28 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX230
+ bl_230 br_230 bl_out_28 br_out_28 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX231
+ bl_231 br_231 bl_out_28 br_out_28 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX232
+ bl_232 br_232 bl_out_29 br_out_29 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX233
+ bl_233 br_233 bl_out_29 br_out_29 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX234
+ bl_234 br_234 bl_out_29 br_out_29 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX235
+ bl_235 br_235 bl_out_29 br_out_29 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX236
+ bl_236 br_236 bl_out_29 br_out_29 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX237
+ bl_237 br_237 bl_out_29 br_out_29 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX238
+ bl_238 br_238 bl_out_29 br_out_29 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX239
+ bl_239 br_239 bl_out_29 br_out_29 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX240
+ bl_240 br_240 bl_out_30 br_out_30 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX241
+ bl_241 br_241 bl_out_30 br_out_30 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX242
+ bl_242 br_242 bl_out_30 br_out_30 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX243
+ bl_243 br_243 bl_out_30 br_out_30 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX244
+ bl_244 br_244 bl_out_30 br_out_30 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX245
+ bl_245 br_245 bl_out_30 br_out_30 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX246
+ bl_246 br_246 bl_out_30 br_out_30 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX247
+ bl_247 br_247 bl_out_30 br_out_30 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX248
+ bl_248 br_248 bl_out_31 br_out_31 sel_0 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX249
+ bl_249 br_249 bl_out_31 br_out_31 sel_1 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX250
+ bl_250 br_250 bl_out_31 br_out_31 sel_2 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX251
+ bl_251 br_251 bl_out_31 br_out_31 sel_3 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX252
+ bl_252 br_252 bl_out_31 br_out_31 sel_4 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX253
+ bl_253 br_253 bl_out_31 br_out_31 sel_5 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX254
+ bl_254 br_254 bl_out_31 br_out_31 sel_6 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
XXMUX255
+ bl_255 br_255 bl_out_31 br_out_31 sel_7 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux
.ENDS sram_1rw0r0w_32_1024_freepdk45_column_mux_array

.SUBCKT write_driver din bl br en vdd gnd
*inverters for enable and data input
minP bl_bar din vdd vdd pmos_vtg w=360.000000n l=50.000000n
minN bl_bar din gnd gnd nmos_vtg w=180.000000n l=50.000000n
moutP en_bar en vdd vdd pmos_vtg w=360.000000n l=50.000000n
moutN en_bar en gnd gnd nmos_vtg w=180.000000n l=50.000000n

*tristate for BL
mout0P int1 bl_bar vdd vdd pmos_vtg w=360.000000n l=50.000000n
mout0P2 bl en_bar int1 vdd pmos_vtg w=360.000000n l=50.000000n
mout0N bl en int2 gnd nmos_vtg w=180.000000n l=50.000000n
mout0N2 int2 bl_bar gnd gnd nmos_vtg w=180.000000n l=50.000000n

*tristate for BR
mout1P int3 din vdd vdd pmos_vtg w=360.000000n l=50.000000n
mout1P2 br en_bar int3 vdd pmos_vtg w=360.000000n l=50.000000n
mout1N br en int4 gnd nmos_vtg w=180.000000n l=50.000000n
mout1N2 int4 din gnd gnd nmos_vtg w=180.000000n l=50.000000n
.ENDS write_driver


.SUBCKT sram_1rw0r0w_32_1024_freepdk45_write_driver_array
+ data_0 data_1 data_2 data_3 data_4 data_5 data_6 data_7 data_8 data_9
+ data_10 data_11 data_12 data_13 data_14 data_15 data_16 data_17
+ data_18 data_19 data_20 data_21 data_22 data_23 data_24 data_25
+ data_26 data_27 data_28 data_29 data_30 data_31 bl_0 br_0 bl_1 br_1
+ bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8
+ bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14
+ bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20
+ br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25
+ bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31
+ br_31 en vdd gnd
* INPUT : data_0 
* INPUT : data_1 
* INPUT : data_2 
* INPUT : data_3 
* INPUT : data_4 
* INPUT : data_5 
* INPUT : data_6 
* INPUT : data_7 
* INPUT : data_8 
* INPUT : data_9 
* INPUT : data_10 
* INPUT : data_11 
* INPUT : data_12 
* INPUT : data_13 
* INPUT : data_14 
* INPUT : data_15 
* INPUT : data_16 
* INPUT : data_17 
* INPUT : data_18 
* INPUT : data_19 
* INPUT : data_20 
* INPUT : data_21 
* INPUT : data_22 
* INPUT : data_23 
* INPUT : data_24 
* INPUT : data_25 
* INPUT : data_26 
* INPUT : data_27 
* INPUT : data_28 
* INPUT : data_29 
* INPUT : data_30 
* INPUT : data_31 
* OUTPUT: bl_0 
* OUTPUT: br_0 
* OUTPUT: bl_1 
* OUTPUT: br_1 
* OUTPUT: bl_2 
* OUTPUT: br_2 
* OUTPUT: bl_3 
* OUTPUT: br_3 
* OUTPUT: bl_4 
* OUTPUT: br_4 
* OUTPUT: bl_5 
* OUTPUT: br_5 
* OUTPUT: bl_6 
* OUTPUT: br_6 
* OUTPUT: bl_7 
* OUTPUT: br_7 
* OUTPUT: bl_8 
* OUTPUT: br_8 
* OUTPUT: bl_9 
* OUTPUT: br_9 
* OUTPUT: bl_10 
* OUTPUT: br_10 
* OUTPUT: bl_11 
* OUTPUT: br_11 
* OUTPUT: bl_12 
* OUTPUT: br_12 
* OUTPUT: bl_13 
* OUTPUT: br_13 
* OUTPUT: bl_14 
* OUTPUT: br_14 
* OUTPUT: bl_15 
* OUTPUT: br_15 
* OUTPUT: bl_16 
* OUTPUT: br_16 
* OUTPUT: bl_17 
* OUTPUT: br_17 
* OUTPUT: bl_18 
* OUTPUT: br_18 
* OUTPUT: bl_19 
* OUTPUT: br_19 
* OUTPUT: bl_20 
* OUTPUT: br_20 
* OUTPUT: bl_21 
* OUTPUT: br_21 
* OUTPUT: bl_22 
* OUTPUT: br_22 
* OUTPUT: bl_23 
* OUTPUT: br_23 
* OUTPUT: bl_24 
* OUTPUT: br_24 
* OUTPUT: bl_25 
* OUTPUT: br_25 
* OUTPUT: bl_26 
* OUTPUT: br_26 
* OUTPUT: bl_27 
* OUTPUT: br_27 
* OUTPUT: bl_28 
* OUTPUT: br_28 
* OUTPUT: bl_29 
* OUTPUT: br_29 
* OUTPUT: bl_30 
* OUTPUT: br_30 
* OUTPUT: bl_31 
* OUTPUT: br_31 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* columns: 256
* word_size 32
Xwrite_driver0
+ data_0 bl_0 br_0 en vdd gnd
+ write_driver
Xwrite_driver8
+ data_1 bl_1 br_1 en vdd gnd
+ write_driver
Xwrite_driver16
+ data_2 bl_2 br_2 en vdd gnd
+ write_driver
Xwrite_driver24
+ data_3 bl_3 br_3 en vdd gnd
+ write_driver
Xwrite_driver32
+ data_4 bl_4 br_4 en vdd gnd
+ write_driver
Xwrite_driver40
+ data_5 bl_5 br_5 en vdd gnd
+ write_driver
Xwrite_driver48
+ data_6 bl_6 br_6 en vdd gnd
+ write_driver
Xwrite_driver56
+ data_7 bl_7 br_7 en vdd gnd
+ write_driver
Xwrite_driver64
+ data_8 bl_8 br_8 en vdd gnd
+ write_driver
Xwrite_driver72
+ data_9 bl_9 br_9 en vdd gnd
+ write_driver
Xwrite_driver80
+ data_10 bl_10 br_10 en vdd gnd
+ write_driver
Xwrite_driver88
+ data_11 bl_11 br_11 en vdd gnd
+ write_driver
Xwrite_driver96
+ data_12 bl_12 br_12 en vdd gnd
+ write_driver
Xwrite_driver104
+ data_13 bl_13 br_13 en vdd gnd
+ write_driver
Xwrite_driver112
+ data_14 bl_14 br_14 en vdd gnd
+ write_driver
Xwrite_driver120
+ data_15 bl_15 br_15 en vdd gnd
+ write_driver
Xwrite_driver128
+ data_16 bl_16 br_16 en vdd gnd
+ write_driver
Xwrite_driver136
+ data_17 bl_17 br_17 en vdd gnd
+ write_driver
Xwrite_driver144
+ data_18 bl_18 br_18 en vdd gnd
+ write_driver
Xwrite_driver152
+ data_19 bl_19 br_19 en vdd gnd
+ write_driver
Xwrite_driver160
+ data_20 bl_20 br_20 en vdd gnd
+ write_driver
Xwrite_driver168
+ data_21 bl_21 br_21 en vdd gnd
+ write_driver
Xwrite_driver176
+ data_22 bl_22 br_22 en vdd gnd
+ write_driver
Xwrite_driver184
+ data_23 bl_23 br_23 en vdd gnd
+ write_driver
Xwrite_driver192
+ data_24 bl_24 br_24 en vdd gnd
+ write_driver
Xwrite_driver200
+ data_25 bl_25 br_25 en vdd gnd
+ write_driver
Xwrite_driver208
+ data_26 bl_26 br_26 en vdd gnd
+ write_driver
Xwrite_driver216
+ data_27 bl_27 br_27 en vdd gnd
+ write_driver
Xwrite_driver224
+ data_28 bl_28 br_28 en vdd gnd
+ write_driver
Xwrite_driver232
+ data_29 bl_29 br_29 en vdd gnd
+ write_driver
Xwrite_driver240
+ data_30 bl_30 br_30 en vdd gnd
+ write_driver
Xwrite_driver248
+ data_31 bl_31 br_31 en vdd gnd
+ write_driver
.ENDS sram_1rw0r0w_32_1024_freepdk45_write_driver_array

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_port_data
+ rbl_bl rbl_br bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5
+ br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11
+ bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17
+ br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22
+ bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28
+ br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33
+ bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39
+ br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44
+ bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50
+ br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55
+ bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61
+ br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66
+ bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72
+ br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77
+ bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83
+ br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88
+ bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94
+ br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99
+ bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104
+ bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109
+ bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114
+ bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119
+ bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124
+ bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129
+ bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134
+ bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139
+ bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144
+ bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149
+ bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154
+ bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159
+ bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164
+ bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169
+ bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174
+ bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179
+ bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184
+ bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189
+ bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194
+ bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199
+ bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204
+ bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209
+ bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214
+ bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219
+ bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224
+ bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229
+ bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234
+ bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239
+ bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244
+ bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249
+ bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254
+ bl_255 br_255 dout_0 dout_1 dout_2 dout_3 dout_4 dout_5 dout_6 dout_7
+ dout_8 dout_9 dout_10 dout_11 dout_12 dout_13 dout_14 dout_15 dout_16
+ dout_17 dout_18 dout_19 dout_20 dout_21 dout_22 dout_23 dout_24
+ dout_25 dout_26 dout_27 dout_28 dout_29 dout_30 dout_31 din_0 din_1
+ din_2 din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10 din_11 din_12
+ din_13 din_14 din_15 din_16 din_17 din_18 din_19 din_20 din_21 din_22
+ din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30 din_31 sel_0
+ sel_1 sel_2 sel_3 sel_4 sel_5 sel_6 sel_7 s_en p_en_bar w_en vdd gnd
* INOUT : rbl_bl 
* INOUT : rbl_br 
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : bl_64 
* INOUT : br_64 
* INOUT : bl_65 
* INOUT : br_65 
* INOUT : bl_66 
* INOUT : br_66 
* INOUT : bl_67 
* INOUT : br_67 
* INOUT : bl_68 
* INOUT : br_68 
* INOUT : bl_69 
* INOUT : br_69 
* INOUT : bl_70 
* INOUT : br_70 
* INOUT : bl_71 
* INOUT : br_71 
* INOUT : bl_72 
* INOUT : br_72 
* INOUT : bl_73 
* INOUT : br_73 
* INOUT : bl_74 
* INOUT : br_74 
* INOUT : bl_75 
* INOUT : br_75 
* INOUT : bl_76 
* INOUT : br_76 
* INOUT : bl_77 
* INOUT : br_77 
* INOUT : bl_78 
* INOUT : br_78 
* INOUT : bl_79 
* INOUT : br_79 
* INOUT : bl_80 
* INOUT : br_80 
* INOUT : bl_81 
* INOUT : br_81 
* INOUT : bl_82 
* INOUT : br_82 
* INOUT : bl_83 
* INOUT : br_83 
* INOUT : bl_84 
* INOUT : br_84 
* INOUT : bl_85 
* INOUT : br_85 
* INOUT : bl_86 
* INOUT : br_86 
* INOUT : bl_87 
* INOUT : br_87 
* INOUT : bl_88 
* INOUT : br_88 
* INOUT : bl_89 
* INOUT : br_89 
* INOUT : bl_90 
* INOUT : br_90 
* INOUT : bl_91 
* INOUT : br_91 
* INOUT : bl_92 
* INOUT : br_92 
* INOUT : bl_93 
* INOUT : br_93 
* INOUT : bl_94 
* INOUT : br_94 
* INOUT : bl_95 
* INOUT : br_95 
* INOUT : bl_96 
* INOUT : br_96 
* INOUT : bl_97 
* INOUT : br_97 
* INOUT : bl_98 
* INOUT : br_98 
* INOUT : bl_99 
* INOUT : br_99 
* INOUT : bl_100 
* INOUT : br_100 
* INOUT : bl_101 
* INOUT : br_101 
* INOUT : bl_102 
* INOUT : br_102 
* INOUT : bl_103 
* INOUT : br_103 
* INOUT : bl_104 
* INOUT : br_104 
* INOUT : bl_105 
* INOUT : br_105 
* INOUT : bl_106 
* INOUT : br_106 
* INOUT : bl_107 
* INOUT : br_107 
* INOUT : bl_108 
* INOUT : br_108 
* INOUT : bl_109 
* INOUT : br_109 
* INOUT : bl_110 
* INOUT : br_110 
* INOUT : bl_111 
* INOUT : br_111 
* INOUT : bl_112 
* INOUT : br_112 
* INOUT : bl_113 
* INOUT : br_113 
* INOUT : bl_114 
* INOUT : br_114 
* INOUT : bl_115 
* INOUT : br_115 
* INOUT : bl_116 
* INOUT : br_116 
* INOUT : bl_117 
* INOUT : br_117 
* INOUT : bl_118 
* INOUT : br_118 
* INOUT : bl_119 
* INOUT : br_119 
* INOUT : bl_120 
* INOUT : br_120 
* INOUT : bl_121 
* INOUT : br_121 
* INOUT : bl_122 
* INOUT : br_122 
* INOUT : bl_123 
* INOUT : br_123 
* INOUT : bl_124 
* INOUT : br_124 
* INOUT : bl_125 
* INOUT : br_125 
* INOUT : bl_126 
* INOUT : br_126 
* INOUT : bl_127 
* INOUT : br_127 
* INOUT : bl_128 
* INOUT : br_128 
* INOUT : bl_129 
* INOUT : br_129 
* INOUT : bl_130 
* INOUT : br_130 
* INOUT : bl_131 
* INOUT : br_131 
* INOUT : bl_132 
* INOUT : br_132 
* INOUT : bl_133 
* INOUT : br_133 
* INOUT : bl_134 
* INOUT : br_134 
* INOUT : bl_135 
* INOUT : br_135 
* INOUT : bl_136 
* INOUT : br_136 
* INOUT : bl_137 
* INOUT : br_137 
* INOUT : bl_138 
* INOUT : br_138 
* INOUT : bl_139 
* INOUT : br_139 
* INOUT : bl_140 
* INOUT : br_140 
* INOUT : bl_141 
* INOUT : br_141 
* INOUT : bl_142 
* INOUT : br_142 
* INOUT : bl_143 
* INOUT : br_143 
* INOUT : bl_144 
* INOUT : br_144 
* INOUT : bl_145 
* INOUT : br_145 
* INOUT : bl_146 
* INOUT : br_146 
* INOUT : bl_147 
* INOUT : br_147 
* INOUT : bl_148 
* INOUT : br_148 
* INOUT : bl_149 
* INOUT : br_149 
* INOUT : bl_150 
* INOUT : br_150 
* INOUT : bl_151 
* INOUT : br_151 
* INOUT : bl_152 
* INOUT : br_152 
* INOUT : bl_153 
* INOUT : br_153 
* INOUT : bl_154 
* INOUT : br_154 
* INOUT : bl_155 
* INOUT : br_155 
* INOUT : bl_156 
* INOUT : br_156 
* INOUT : bl_157 
* INOUT : br_157 
* INOUT : bl_158 
* INOUT : br_158 
* INOUT : bl_159 
* INOUT : br_159 
* INOUT : bl_160 
* INOUT : br_160 
* INOUT : bl_161 
* INOUT : br_161 
* INOUT : bl_162 
* INOUT : br_162 
* INOUT : bl_163 
* INOUT : br_163 
* INOUT : bl_164 
* INOUT : br_164 
* INOUT : bl_165 
* INOUT : br_165 
* INOUT : bl_166 
* INOUT : br_166 
* INOUT : bl_167 
* INOUT : br_167 
* INOUT : bl_168 
* INOUT : br_168 
* INOUT : bl_169 
* INOUT : br_169 
* INOUT : bl_170 
* INOUT : br_170 
* INOUT : bl_171 
* INOUT : br_171 
* INOUT : bl_172 
* INOUT : br_172 
* INOUT : bl_173 
* INOUT : br_173 
* INOUT : bl_174 
* INOUT : br_174 
* INOUT : bl_175 
* INOUT : br_175 
* INOUT : bl_176 
* INOUT : br_176 
* INOUT : bl_177 
* INOUT : br_177 
* INOUT : bl_178 
* INOUT : br_178 
* INOUT : bl_179 
* INOUT : br_179 
* INOUT : bl_180 
* INOUT : br_180 
* INOUT : bl_181 
* INOUT : br_181 
* INOUT : bl_182 
* INOUT : br_182 
* INOUT : bl_183 
* INOUT : br_183 
* INOUT : bl_184 
* INOUT : br_184 
* INOUT : bl_185 
* INOUT : br_185 
* INOUT : bl_186 
* INOUT : br_186 
* INOUT : bl_187 
* INOUT : br_187 
* INOUT : bl_188 
* INOUT : br_188 
* INOUT : bl_189 
* INOUT : br_189 
* INOUT : bl_190 
* INOUT : br_190 
* INOUT : bl_191 
* INOUT : br_191 
* INOUT : bl_192 
* INOUT : br_192 
* INOUT : bl_193 
* INOUT : br_193 
* INOUT : bl_194 
* INOUT : br_194 
* INOUT : bl_195 
* INOUT : br_195 
* INOUT : bl_196 
* INOUT : br_196 
* INOUT : bl_197 
* INOUT : br_197 
* INOUT : bl_198 
* INOUT : br_198 
* INOUT : bl_199 
* INOUT : br_199 
* INOUT : bl_200 
* INOUT : br_200 
* INOUT : bl_201 
* INOUT : br_201 
* INOUT : bl_202 
* INOUT : br_202 
* INOUT : bl_203 
* INOUT : br_203 
* INOUT : bl_204 
* INOUT : br_204 
* INOUT : bl_205 
* INOUT : br_205 
* INOUT : bl_206 
* INOUT : br_206 
* INOUT : bl_207 
* INOUT : br_207 
* INOUT : bl_208 
* INOUT : br_208 
* INOUT : bl_209 
* INOUT : br_209 
* INOUT : bl_210 
* INOUT : br_210 
* INOUT : bl_211 
* INOUT : br_211 
* INOUT : bl_212 
* INOUT : br_212 
* INOUT : bl_213 
* INOUT : br_213 
* INOUT : bl_214 
* INOUT : br_214 
* INOUT : bl_215 
* INOUT : br_215 
* INOUT : bl_216 
* INOUT : br_216 
* INOUT : bl_217 
* INOUT : br_217 
* INOUT : bl_218 
* INOUT : br_218 
* INOUT : bl_219 
* INOUT : br_219 
* INOUT : bl_220 
* INOUT : br_220 
* INOUT : bl_221 
* INOUT : br_221 
* INOUT : bl_222 
* INOUT : br_222 
* INOUT : bl_223 
* INOUT : br_223 
* INOUT : bl_224 
* INOUT : br_224 
* INOUT : bl_225 
* INOUT : br_225 
* INOUT : bl_226 
* INOUT : br_226 
* INOUT : bl_227 
* INOUT : br_227 
* INOUT : bl_228 
* INOUT : br_228 
* INOUT : bl_229 
* INOUT : br_229 
* INOUT : bl_230 
* INOUT : br_230 
* INOUT : bl_231 
* INOUT : br_231 
* INOUT : bl_232 
* INOUT : br_232 
* INOUT : bl_233 
* INOUT : br_233 
* INOUT : bl_234 
* INOUT : br_234 
* INOUT : bl_235 
* INOUT : br_235 
* INOUT : bl_236 
* INOUT : br_236 
* INOUT : bl_237 
* INOUT : br_237 
* INOUT : bl_238 
* INOUT : br_238 
* INOUT : bl_239 
* INOUT : br_239 
* INOUT : bl_240 
* INOUT : br_240 
* INOUT : bl_241 
* INOUT : br_241 
* INOUT : bl_242 
* INOUT : br_242 
* INOUT : bl_243 
* INOUT : br_243 
* INOUT : bl_244 
* INOUT : br_244 
* INOUT : bl_245 
* INOUT : br_245 
* INOUT : bl_246 
* INOUT : br_246 
* INOUT : bl_247 
* INOUT : br_247 
* INOUT : bl_248 
* INOUT : br_248 
* INOUT : bl_249 
* INOUT : br_249 
* INOUT : bl_250 
* INOUT : br_250 
* INOUT : bl_251 
* INOUT : br_251 
* INOUT : bl_252 
* INOUT : br_252 
* INOUT : bl_253 
* INOUT : br_253 
* INOUT : bl_254 
* INOUT : br_254 
* INOUT : bl_255 
* INOUT : br_255 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* OUTPUT: dout_7 
* OUTPUT: dout_8 
* OUTPUT: dout_9 
* OUTPUT: dout_10 
* OUTPUT: dout_11 
* OUTPUT: dout_12 
* OUTPUT: dout_13 
* OUTPUT: dout_14 
* OUTPUT: dout_15 
* OUTPUT: dout_16 
* OUTPUT: dout_17 
* OUTPUT: dout_18 
* OUTPUT: dout_19 
* OUTPUT: dout_20 
* OUTPUT: dout_21 
* OUTPUT: dout_22 
* OUTPUT: dout_23 
* OUTPUT: dout_24 
* OUTPUT: dout_25 
* OUTPUT: dout_26 
* OUTPUT: dout_27 
* OUTPUT: dout_28 
* OUTPUT: dout_29 
* OUTPUT: dout_30 
* OUTPUT: dout_31 
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* INPUT : din_7 
* INPUT : din_8 
* INPUT : din_9 
* INPUT : din_10 
* INPUT : din_11 
* INPUT : din_12 
* INPUT : din_13 
* INPUT : din_14 
* INPUT : din_15 
* INPUT : din_16 
* INPUT : din_17 
* INPUT : din_18 
* INPUT : din_19 
* INPUT : din_20 
* INPUT : din_21 
* INPUT : din_22 
* INPUT : din_23 
* INPUT : din_24 
* INPUT : din_25 
* INPUT : din_26 
* INPUT : din_27 
* INPUT : din_28 
* INPUT : din_29 
* INPUT : din_30 
* INPUT : din_31 
* INPUT : sel_0 
* INPUT : sel_1 
* INPUT : sel_2 
* INPUT : sel_3 
* INPUT : sel_4 
* INPUT : sel_5 
* INPUT : sel_6 
* INPUT : sel_7 
* INPUT : s_en 
* INPUT : p_en_bar 
* INPUT : w_en 
* POWER : vdd 
* GROUND: gnd 
Xprecharge_array0
+ rbl_bl rbl_br bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5
+ br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11
+ bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17
+ br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22
+ bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28
+ br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33
+ bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39
+ br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44
+ bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50
+ br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55
+ bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61
+ br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66
+ bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72
+ br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77
+ bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83
+ br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88
+ bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94
+ br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99
+ bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104
+ bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109
+ bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114
+ bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119
+ bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124
+ bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129
+ bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134
+ bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139
+ bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144
+ bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149
+ bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154
+ bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159
+ bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164
+ bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169
+ bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174
+ bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179
+ bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184
+ bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189
+ bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194
+ bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199
+ bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204
+ bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209
+ bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214
+ bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219
+ bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224
+ bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229
+ bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234
+ bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239
+ bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244
+ bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249
+ bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254
+ bl_255 br_255 p_en_bar vdd
+ sram_1rw0r0w_32_1024_freepdk45_precharge_array
Xsense_amp_array0
+ dout_0 bl_out_0 br_out_0 dout_1 bl_out_1 br_out_1 dout_2 bl_out_2
+ br_out_2 dout_3 bl_out_3 br_out_3 dout_4 bl_out_4 br_out_4 dout_5
+ bl_out_5 br_out_5 dout_6 bl_out_6 br_out_6 dout_7 bl_out_7 br_out_7
+ dout_8 bl_out_8 br_out_8 dout_9 bl_out_9 br_out_9 dout_10 bl_out_10
+ br_out_10 dout_11 bl_out_11 br_out_11 dout_12 bl_out_12 br_out_12
+ dout_13 bl_out_13 br_out_13 dout_14 bl_out_14 br_out_14 dout_15
+ bl_out_15 br_out_15 dout_16 bl_out_16 br_out_16 dout_17 bl_out_17
+ br_out_17 dout_18 bl_out_18 br_out_18 dout_19 bl_out_19 br_out_19
+ dout_20 bl_out_20 br_out_20 dout_21 bl_out_21 br_out_21 dout_22
+ bl_out_22 br_out_22 dout_23 bl_out_23 br_out_23 dout_24 bl_out_24
+ br_out_24 dout_25 bl_out_25 br_out_25 dout_26 bl_out_26 br_out_26
+ dout_27 bl_out_27 br_out_27 dout_28 bl_out_28 br_out_28 dout_29
+ bl_out_29 br_out_29 dout_30 bl_out_30 br_out_30 dout_31 bl_out_31
+ br_out_31 s_en vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_sense_amp_array
Xwrite_driver_array0
+ din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10
+ din_11 din_12 din_13 din_14 din_15 din_16 din_17 din_18 din_19 din_20
+ din_21 din_22 din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30
+ din_31 bl_out_0 br_out_0 bl_out_1 br_out_1 bl_out_2 br_out_2 bl_out_3
+ br_out_3 bl_out_4 br_out_4 bl_out_5 br_out_5 bl_out_6 br_out_6
+ bl_out_7 br_out_7 bl_out_8 br_out_8 bl_out_9 br_out_9 bl_out_10
+ br_out_10 bl_out_11 br_out_11 bl_out_12 br_out_12 bl_out_13 br_out_13
+ bl_out_14 br_out_14 bl_out_15 br_out_15 bl_out_16 br_out_16 bl_out_17
+ br_out_17 bl_out_18 br_out_18 bl_out_19 br_out_19 bl_out_20 br_out_20
+ bl_out_21 br_out_21 bl_out_22 br_out_22 bl_out_23 br_out_23 bl_out_24
+ br_out_24 bl_out_25 br_out_25 bl_out_26 br_out_26 bl_out_27 br_out_27
+ bl_out_28 br_out_28 bl_out_29 br_out_29 bl_out_30 br_out_30 bl_out_31
+ br_out_31 w_en vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_write_driver_array
Xcolumn_mux_array0
+ bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6
+ bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12
+ bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18
+ br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23
+ bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29
+ br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34
+ bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40
+ br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45
+ bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51
+ br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56
+ bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62
+ br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67
+ bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73
+ br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78
+ bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84
+ br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89
+ bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95
+ br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100
+ bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105
+ bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110
+ bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115
+ bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120
+ bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125
+ bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130
+ bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135
+ bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140
+ bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145
+ bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150
+ bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155
+ bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160
+ bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165
+ bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170
+ bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175
+ bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180
+ bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185
+ bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190
+ bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195
+ bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200
+ bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205
+ bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210
+ bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215
+ bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220
+ bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225
+ bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230
+ bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235
+ bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240
+ bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245
+ bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250
+ bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255
+ sel_0 sel_1 sel_2 sel_3 sel_4 sel_5 sel_6 sel_7 bl_out_0 br_out_0
+ bl_out_1 br_out_1 bl_out_2 br_out_2 bl_out_3 br_out_3 bl_out_4
+ br_out_4 bl_out_5 br_out_5 bl_out_6 br_out_6 bl_out_7 br_out_7
+ bl_out_8 br_out_8 bl_out_9 br_out_9 bl_out_10 br_out_10 bl_out_11
+ br_out_11 bl_out_12 br_out_12 bl_out_13 br_out_13 bl_out_14 br_out_14
+ bl_out_15 br_out_15 bl_out_16 br_out_16 bl_out_17 br_out_17 bl_out_18
+ br_out_18 bl_out_19 br_out_19 bl_out_20 br_out_20 bl_out_21 br_out_21
+ bl_out_22 br_out_22 bl_out_23 br_out_23 bl_out_24 br_out_24 bl_out_25
+ br_out_25 bl_out_26 br_out_26 bl_out_27 br_out_27 bl_out_28 br_out_28
+ bl_out_29 br_out_29 bl_out_30 br_out_30 bl_out_31 br_out_31 gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_mux_array
.ENDS sram_1rw0r0w_32_1024_freepdk45_port_data

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_bank
+ dout0_0 dout0_1 dout0_2 dout0_3 dout0_4 dout0_5 dout0_6 dout0_7
+ dout0_8 dout0_9 dout0_10 dout0_11 dout0_12 dout0_13 dout0_14 dout0_15
+ dout0_16 dout0_17 dout0_18 dout0_19 dout0_20 dout0_21 dout0_22
+ dout0_23 dout0_24 dout0_25 dout0_26 dout0_27 dout0_28 dout0_29
+ dout0_30 dout0_31 rbl_bl_0_0 din0_0 din0_1 din0_2 din0_3 din0_4 din0_5
+ din0_6 din0_7 din0_8 din0_9 din0_10 din0_11 din0_12 din0_13 din0_14
+ din0_15 din0_16 din0_17 din0_18 din0_19 din0_20 din0_21 din0_22
+ din0_23 din0_24 din0_25 din0_26 din0_27 din0_28 din0_29 din0_30
+ din0_31 addr0_0 addr0_1 addr0_2 addr0_3 addr0_4 addr0_5 addr0_6
+ addr0_7 addr0_8 addr0_9 s_en0 p_en_bar0 w_en0 wl_en0 vdd gnd
* OUTPUT: dout0_0 
* OUTPUT: dout0_1 
* OUTPUT: dout0_2 
* OUTPUT: dout0_3 
* OUTPUT: dout0_4 
* OUTPUT: dout0_5 
* OUTPUT: dout0_6 
* OUTPUT: dout0_7 
* OUTPUT: dout0_8 
* OUTPUT: dout0_9 
* OUTPUT: dout0_10 
* OUTPUT: dout0_11 
* OUTPUT: dout0_12 
* OUTPUT: dout0_13 
* OUTPUT: dout0_14 
* OUTPUT: dout0_15 
* OUTPUT: dout0_16 
* OUTPUT: dout0_17 
* OUTPUT: dout0_18 
* OUTPUT: dout0_19 
* OUTPUT: dout0_20 
* OUTPUT: dout0_21 
* OUTPUT: dout0_22 
* OUTPUT: dout0_23 
* OUTPUT: dout0_24 
* OUTPUT: dout0_25 
* OUTPUT: dout0_26 
* OUTPUT: dout0_27 
* OUTPUT: dout0_28 
* OUTPUT: dout0_29 
* OUTPUT: dout0_30 
* OUTPUT: dout0_31 
* OUTPUT: rbl_bl_0_0 
* INPUT : din0_0 
* INPUT : din0_1 
* INPUT : din0_2 
* INPUT : din0_3 
* INPUT : din0_4 
* INPUT : din0_5 
* INPUT : din0_6 
* INPUT : din0_7 
* INPUT : din0_8 
* INPUT : din0_9 
* INPUT : din0_10 
* INPUT : din0_11 
* INPUT : din0_12 
* INPUT : din0_13 
* INPUT : din0_14 
* INPUT : din0_15 
* INPUT : din0_16 
* INPUT : din0_17 
* INPUT : din0_18 
* INPUT : din0_19 
* INPUT : din0_20 
* INPUT : din0_21 
* INPUT : din0_22 
* INPUT : din0_23 
* INPUT : din0_24 
* INPUT : din0_25 
* INPUT : din0_26 
* INPUT : din0_27 
* INPUT : din0_28 
* INPUT : din0_29 
* INPUT : din0_30 
* INPUT : din0_31 
* INPUT : addr0_0 
* INPUT : addr0_1 
* INPUT : addr0_2 
* INPUT : addr0_3 
* INPUT : addr0_4 
* INPUT : addr0_5 
* INPUT : addr0_6 
* INPUT : addr0_7 
* INPUT : addr0_8 
* INPUT : addr0_9 
* INPUT : s_en0 
* INPUT : p_en_bar0 
* INPUT : w_en0 
* INPUT : wl_en0 
* POWER : vdd 
* GROUND: gnd 
Xbitcell_array
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64
+ bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68
+ bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72
+ bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76
+ bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80
+ bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84
+ bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88
+ bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92
+ bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96
+ bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100
+ bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104
+ br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107
+ bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111
+ br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114
+ bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118
+ br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121
+ bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125
+ br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128
+ bl_0_129 br_0_129 bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132
+ br_0_132 bl_0_133 br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135
+ bl_0_136 br_0_136 bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139
+ br_0_139 bl_0_140 br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142
+ bl_0_143 br_0_143 bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146
+ br_0_146 bl_0_147 br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149
+ bl_0_150 br_0_150 bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153
+ br_0_153 bl_0_154 br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156
+ bl_0_157 br_0_157 bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160
+ br_0_160 bl_0_161 br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163
+ bl_0_164 br_0_164 bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167
+ br_0_167 bl_0_168 br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170
+ bl_0_171 br_0_171 bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174
+ br_0_174 bl_0_175 br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177
+ bl_0_178 br_0_178 bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181
+ br_0_181 bl_0_182 br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184
+ bl_0_185 br_0_185 bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188
+ br_0_188 bl_0_189 br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191
+ bl_0_192 br_0_192 bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195
+ br_0_195 bl_0_196 br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198
+ bl_0_199 br_0_199 bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202
+ br_0_202 bl_0_203 br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205
+ bl_0_206 br_0_206 bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209
+ br_0_209 bl_0_210 br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212
+ bl_0_213 br_0_213 bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216
+ br_0_216 bl_0_217 br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219
+ bl_0_220 br_0_220 bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223
+ br_0_223 bl_0_224 br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226
+ bl_0_227 br_0_227 bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230
+ br_0_230 bl_0_231 br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233
+ bl_0_234 br_0_234 bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237
+ br_0_237 bl_0_238 br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240
+ bl_0_241 br_0_241 bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244
+ br_0_244 bl_0_245 br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247
+ bl_0_248 br_0_248 bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251
+ br_0_251 bl_0_252 br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254
+ bl_0_255 br_0_255 rbl_wl0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5
+ wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14
+ wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22
+ wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30
+ wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38
+ wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46
+ wl_0_47 wl_0_48 wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54
+ wl_0_55 wl_0_56 wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62
+ wl_0_63 wl_0_64 wl_0_65 wl_0_66 wl_0_67 wl_0_68 wl_0_69 wl_0_70
+ wl_0_71 wl_0_72 wl_0_73 wl_0_74 wl_0_75 wl_0_76 wl_0_77 wl_0_78
+ wl_0_79 wl_0_80 wl_0_81 wl_0_82 wl_0_83 wl_0_84 wl_0_85 wl_0_86
+ wl_0_87 wl_0_88 wl_0_89 wl_0_90 wl_0_91 wl_0_92 wl_0_93 wl_0_94
+ wl_0_95 wl_0_96 wl_0_97 wl_0_98 wl_0_99 wl_0_100 wl_0_101 wl_0_102
+ wl_0_103 wl_0_104 wl_0_105 wl_0_106 wl_0_107 wl_0_108 wl_0_109
+ wl_0_110 wl_0_111 wl_0_112 wl_0_113 wl_0_114 wl_0_115 wl_0_116
+ wl_0_117 wl_0_118 wl_0_119 wl_0_120 wl_0_121 wl_0_122 wl_0_123
+ wl_0_124 wl_0_125 wl_0_126 wl_0_127 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_capped_replica_bitcell_array
Xport_data0
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64
+ bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68
+ bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72
+ bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76
+ bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80
+ bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84
+ bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88
+ bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92
+ bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96
+ bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100
+ bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104
+ br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107
+ bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111
+ br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114
+ bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118
+ br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121
+ bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125
+ br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128
+ bl_0_129 br_0_129 bl_0_130 br_0_130 bl_0_131 br_0_131 bl_0_132
+ br_0_132 bl_0_133 br_0_133 bl_0_134 br_0_134 bl_0_135 br_0_135
+ bl_0_136 br_0_136 bl_0_137 br_0_137 bl_0_138 br_0_138 bl_0_139
+ br_0_139 bl_0_140 br_0_140 bl_0_141 br_0_141 bl_0_142 br_0_142
+ bl_0_143 br_0_143 bl_0_144 br_0_144 bl_0_145 br_0_145 bl_0_146
+ br_0_146 bl_0_147 br_0_147 bl_0_148 br_0_148 bl_0_149 br_0_149
+ bl_0_150 br_0_150 bl_0_151 br_0_151 bl_0_152 br_0_152 bl_0_153
+ br_0_153 bl_0_154 br_0_154 bl_0_155 br_0_155 bl_0_156 br_0_156
+ bl_0_157 br_0_157 bl_0_158 br_0_158 bl_0_159 br_0_159 bl_0_160
+ br_0_160 bl_0_161 br_0_161 bl_0_162 br_0_162 bl_0_163 br_0_163
+ bl_0_164 br_0_164 bl_0_165 br_0_165 bl_0_166 br_0_166 bl_0_167
+ br_0_167 bl_0_168 br_0_168 bl_0_169 br_0_169 bl_0_170 br_0_170
+ bl_0_171 br_0_171 bl_0_172 br_0_172 bl_0_173 br_0_173 bl_0_174
+ br_0_174 bl_0_175 br_0_175 bl_0_176 br_0_176 bl_0_177 br_0_177
+ bl_0_178 br_0_178 bl_0_179 br_0_179 bl_0_180 br_0_180 bl_0_181
+ br_0_181 bl_0_182 br_0_182 bl_0_183 br_0_183 bl_0_184 br_0_184
+ bl_0_185 br_0_185 bl_0_186 br_0_186 bl_0_187 br_0_187 bl_0_188
+ br_0_188 bl_0_189 br_0_189 bl_0_190 br_0_190 bl_0_191 br_0_191
+ bl_0_192 br_0_192 bl_0_193 br_0_193 bl_0_194 br_0_194 bl_0_195
+ br_0_195 bl_0_196 br_0_196 bl_0_197 br_0_197 bl_0_198 br_0_198
+ bl_0_199 br_0_199 bl_0_200 br_0_200 bl_0_201 br_0_201 bl_0_202
+ br_0_202 bl_0_203 br_0_203 bl_0_204 br_0_204 bl_0_205 br_0_205
+ bl_0_206 br_0_206 bl_0_207 br_0_207 bl_0_208 br_0_208 bl_0_209
+ br_0_209 bl_0_210 br_0_210 bl_0_211 br_0_211 bl_0_212 br_0_212
+ bl_0_213 br_0_213 bl_0_214 br_0_214 bl_0_215 br_0_215 bl_0_216
+ br_0_216 bl_0_217 br_0_217 bl_0_218 br_0_218 bl_0_219 br_0_219
+ bl_0_220 br_0_220 bl_0_221 br_0_221 bl_0_222 br_0_222 bl_0_223
+ br_0_223 bl_0_224 br_0_224 bl_0_225 br_0_225 bl_0_226 br_0_226
+ bl_0_227 br_0_227 bl_0_228 br_0_228 bl_0_229 br_0_229 bl_0_230
+ br_0_230 bl_0_231 br_0_231 bl_0_232 br_0_232 bl_0_233 br_0_233
+ bl_0_234 br_0_234 bl_0_235 br_0_235 bl_0_236 br_0_236 bl_0_237
+ br_0_237 bl_0_238 br_0_238 bl_0_239 br_0_239 bl_0_240 br_0_240
+ bl_0_241 br_0_241 bl_0_242 br_0_242 bl_0_243 br_0_243 bl_0_244
+ br_0_244 bl_0_245 br_0_245 bl_0_246 br_0_246 bl_0_247 br_0_247
+ bl_0_248 br_0_248 bl_0_249 br_0_249 bl_0_250 br_0_250 bl_0_251
+ br_0_251 bl_0_252 br_0_252 bl_0_253 br_0_253 bl_0_254 br_0_254
+ bl_0_255 br_0_255 dout0_0 dout0_1 dout0_2 dout0_3 dout0_4 dout0_5
+ dout0_6 dout0_7 dout0_8 dout0_9 dout0_10 dout0_11 dout0_12 dout0_13
+ dout0_14 dout0_15 dout0_16 dout0_17 dout0_18 dout0_19 dout0_20
+ dout0_21 dout0_22 dout0_23 dout0_24 dout0_25 dout0_26 dout0_27
+ dout0_28 dout0_29 dout0_30 dout0_31 din0_0 din0_1 din0_2 din0_3 din0_4
+ din0_5 din0_6 din0_7 din0_8 din0_9 din0_10 din0_11 din0_12 din0_13
+ din0_14 din0_15 din0_16 din0_17 din0_18 din0_19 din0_20 din0_21
+ din0_22 din0_23 din0_24 din0_25 din0_26 din0_27 din0_28 din0_29
+ din0_30 din0_31 sel0_0 sel0_1 sel0_2 sel0_3 sel0_4 sel0_5 sel0_6
+ sel0_7 s_en0 p_en_bar0 w_en0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_port_data
Xport_address0
+ addr0_3 addr0_4 addr0_5 addr0_6 addr0_7 addr0_8 addr0_9 wl_en0 wl_0_0
+ wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10
+ wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18
+ wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26
+ wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34
+ wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42
+ wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50
+ wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57 wl_0_58
+ wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 wl_0_65 wl_0_66
+ wl_0_67 wl_0_68 wl_0_69 wl_0_70 wl_0_71 wl_0_72 wl_0_73 wl_0_74
+ wl_0_75 wl_0_76 wl_0_77 wl_0_78 wl_0_79 wl_0_80 wl_0_81 wl_0_82
+ wl_0_83 wl_0_84 wl_0_85 wl_0_86 wl_0_87 wl_0_88 wl_0_89 wl_0_90
+ wl_0_91 wl_0_92 wl_0_93 wl_0_94 wl_0_95 wl_0_96 wl_0_97 wl_0_98
+ wl_0_99 wl_0_100 wl_0_101 wl_0_102 wl_0_103 wl_0_104 wl_0_105 wl_0_106
+ wl_0_107 wl_0_108 wl_0_109 wl_0_110 wl_0_111 wl_0_112 wl_0_113
+ wl_0_114 wl_0_115 wl_0_116 wl_0_117 wl_0_118 wl_0_119 wl_0_120
+ wl_0_121 wl_0_122 wl_0_123 wl_0_124 wl_0_125 wl_0_126 wl_0_127 rbl_wl0
+ vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_port_address
Xcol_address_decoder0
+ addr0_0 addr0_1 addr0_2 sel0_0 sel0_1 sel0_2 sel0_3 sel0_4 sel0_5
+ sel0_6 sel0_7 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_column_decoder
.ENDS sram_1rw0r0w_32_1024_freepdk45_bank

* spice ptx M{0} {1} nmos_vtg m=4 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

* spice ptx M{0} {1} pmos_vtg m=4 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pinv_5
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 12
Mpinv_pmos Z A vdd vdd pmos_vtg m=4 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=4 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pinv_5

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pdriver_0
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [12]
Xbuf_inv1
+ A Z vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_5
.ENDS sram_1rw0r0w_32_1024_freepdk45_pdriver_0

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pnand2_0
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Mpnand2_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_nmos1 Z B net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand2_nmos2 net1 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pnand2_0

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pand2
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 12
Xpand2_nand
+ A B zb_int vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pnand2_0
Xpand2_inv
+ zb_int Z vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pdriver_0
.ENDS sram_1rw0r0w_32_1024_freepdk45_pand2

* spice ptx M{0} {1} nmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

* spice ptx M{0} {1} pmos_vtg m=1 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pinv_8
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 3
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pinv_8

* spice ptx M{0} {1} nmos_vtg m=3 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

* spice ptx M{0} {1} pmos_vtg m=3 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pinv_9
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 9
Mpinv_pmos Z A vdd vdd pmos_vtg m=3 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=3 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pinv_9

* spice ptx M{0} {1} nmos_vtg m=8 w=0.305u l=0.05u pd=0.71u ps=0.71u as=0.04p ad=0.04p

* spice ptx M{0} {1} pmos_vtg m=8 w=0.91u l=0.05u pd=1.92u ps=1.92u as=0.11p ad=0.11p

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pinv_10
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 27
Mpinv_pmos Z A vdd vdd pmos_vtg m=8 w=0.91u l=0.05u pd=1.92u ps=1.92u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=8 w=0.305u l=0.05u pd=0.71u ps=0.71u as=0.04p ad=0.04p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pinv_10

* spice ptx M{0} {1} pmos_vtg m=24 w=0.9u l=0.05u pd=1.90u ps=1.90u as=0.11p ad=0.11p

* spice ptx M{0} {1} nmos_vtg m=24 w=0.3u l=0.05u pd=0.70u ps=0.70u as=0.04p ad=0.04p

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pinv_11
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 80
Mpinv_pmos Z A vdd vdd pmos_vtg m=24 w=0.9u l=0.05u pd=1.90u ps=1.90u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=24 w=0.3u l=0.05u pd=0.70u ps=0.70u as=0.04p ad=0.04p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pinv_11

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pdriver_1
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 3, 9, 27, 80]
Xbuf_inv1
+ A Zb1_int vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_1
Xbuf_inv2
+ Zb1_int Zb2_int vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_1
Xbuf_inv3
+ Zb2_int Zb3_int vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_8
Xbuf_inv4
+ Zb3_int Zb4_int vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_9
Xbuf_inv5
+ Zb4_int Zb5_int vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_10
Xbuf_inv6
+ Zb5_int Z vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_11
.ENDS sram_1rw0r0w_32_1024_freepdk45_pdriver_1

* spice ptx M{0} {1} pmos_vtg m=12 w=0.9u l=0.05u pd=1.90u ps=1.90u as=0.11p ad=0.11p

* spice ptx M{0} {1} nmos_vtg m=12 w=0.3u l=0.05u pd=0.70u ps=0.70u as=0.04p ad=0.04p

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pinv_14
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 40
Mpinv_pmos Z A vdd vdd pmos_vtg m=12 w=0.9u l=0.05u pd=1.90u ps=1.90u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=12 w=0.3u l=0.05u pd=0.70u ps=0.70u as=0.04p ad=0.04p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pinv_14

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pdriver_3
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [40]
Xbuf_inv1
+ A Z vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_14
.ENDS sram_1rw0r0w_32_1024_freepdk45_pdriver_3

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pand3_0
+ A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 40
Xpand3_nand
+ A B C zb_int vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pnand3_0
Xpand3_inv
+ zb_int Z vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pdriver_3
.ENDS sram_1rw0r0w_32_1024_freepdk45_pand3_0

* spice ptx M{0} {1} pmos_vtg m=1 w=0.54u l=0.05u pd=1.18u ps=1.18u as=0.07p ad=0.07p

* spice ptx M{0} {1} nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pinv_3
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 2
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.54u l=0.05u pd=1.18u ps=1.18u as=0.07p ad=0.07p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pinv_3

* spice ptx M{0} {1} pmos_vtg m=2 w=0.54u l=0.05u pd=1.18u ps=1.18u as=0.07p ad=0.07p

* spice ptx M{0} {1} nmos_vtg m=2 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pinv_4
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 4
Mpinv_pmos Z A vdd vdd pmos_vtg m=2 w=0.54u l=0.05u pd=1.18u ps=1.18u as=0.07p ad=0.07p
Mpinv_nmos Z A gnd gnd nmos_vtg m=2 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pinv_4

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_dff_buf_0
+ D Q Qb clk vdd gnd
* INPUT : D 
* OUTPUT: Q 
* OUTPUT: Qb 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* inv1: 2 inv2: 4
Xdff_buf_dff
+ D qint clk vdd gnd
+ dff
Xdff_buf_inv1
+ qint Qb vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_3
Xdff_buf_inv2
+ Qb Q vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_4
.ENDS sram_1rw0r0w_32_1024_freepdk45_dff_buf_0

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_dff_buf_array
+ din_0 din_1 dout_0 dout_bar_0 dout_1 dout_bar_1 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* OUTPUT: dout_0 
* OUTPUT: dout_bar_0 
* OUTPUT: dout_1 
* OUTPUT: dout_bar_1 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 2 cols: 1
* inv1: 2 inv2: 4
Xdff_r0_c0
+ din_0 dout_0 dout_bar_0 clk vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_dff_buf_0
Xdff_r1_c0
+ din_1 dout_1 dout_bar_1 clk vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_dff_buf_0
.ENDS sram_1rw0r0w_32_1024_freepdk45_dff_buf_array

* spice ptx M{0} {1} nmos_vtg m=9 w=0.28u l=0.05u pd=0.66u ps=0.66u as=0.04p ad=0.04p

* spice ptx M{0} {1} pmos_vtg m=9 w=0.84u l=0.05u pd=1.78u ps=1.78u as=0.10p ad=0.10p

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pinv_16
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 28
Mpinv_pmos Z A vdd vdd pmos_vtg m=9 w=0.84u l=0.05u pd=1.78u ps=1.78u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=9 w=0.28u l=0.05u pd=0.66u ps=0.66u as=0.04p ad=0.04p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pinv_16

* spice ptx M{0} {1} nmos_vtg m=25 w=0.305u l=0.05u pd=0.71u ps=0.71u as=0.04p ad=0.04p

* spice ptx M{0} {1} pmos_vtg m=25 w=0.9175u l=0.05u pd=1.94u ps=1.94u as=0.11p ad=0.11p

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pinv_17
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 85
Mpinv_pmos Z A vdd vdd pmos_vtg m=25 w=0.9175u l=0.05u pd=1.94u ps=1.94u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=25 w=0.305u l=0.05u pd=0.71u ps=0.71u as=0.04p ad=0.04p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pinv_17

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pdriver_5
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 3, 9, 28, 85]
Xbuf_inv1
+ A Zb1_int vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_1
Xbuf_inv2
+ Zb1_int Zb2_int vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_1
Xbuf_inv3
+ Zb2_int Zb3_int vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_8
Xbuf_inv4
+ Zb3_int Zb4_int vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_9
Xbuf_inv5
+ Zb4_int Zb5_int vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_16
Xbuf_inv6
+ Zb5_int Z vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_17
.ENDS sram_1rw0r0w_32_1024_freepdk45_pdriver_5

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pinv_18
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pinv_18

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_delay_chain
+ in out vdd gnd
* INPUT : in 
* OUTPUT: out 
* POWER : vdd 
* GROUND: gnd 
* fanouts: [4, 4, 4, 4, 4, 4, 4, 4, 4]
Xdinv0
+ in dout_1 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_0_0
+ dout_1 n_0_0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_0_1
+ dout_1 n_0_1 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_0_2
+ dout_1 n_0_2 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_0_3
+ dout_1 n_0_3 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdinv1
+ dout_1 dout_2 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_1_0
+ dout_2 n_1_0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_1_1
+ dout_2 n_1_1 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_1_2
+ dout_2 n_1_2 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_1_3
+ dout_2 n_1_3 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdinv2
+ dout_2 dout_3 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_2_0
+ dout_3 n_2_0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_2_1
+ dout_3 n_2_1 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_2_2
+ dout_3 n_2_2 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_2_3
+ dout_3 n_2_3 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdinv3
+ dout_3 dout_4 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_3_0
+ dout_4 n_3_0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_3_1
+ dout_4 n_3_1 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_3_2
+ dout_4 n_3_2 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_3_3
+ dout_4 n_3_3 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdinv4
+ dout_4 dout_5 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_4_0
+ dout_5 n_4_0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_4_1
+ dout_5 n_4_1 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_4_2
+ dout_5 n_4_2 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_4_3
+ dout_5 n_4_3 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdinv5
+ dout_5 dout_6 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_5_0
+ dout_6 n_5_0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_5_1
+ dout_6 n_5_1 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_5_2
+ dout_6 n_5_2 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_5_3
+ dout_6 n_5_3 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdinv6
+ dout_6 dout_7 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_6_0
+ dout_7 n_6_0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_6_1
+ dout_7 n_6_1 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_6_2
+ dout_7 n_6_2 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_6_3
+ dout_7 n_6_3 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdinv7
+ dout_7 dout_8 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_7_0
+ dout_8 n_7_0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_7_1
+ dout_8 n_7_1 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_7_2
+ dout_8 n_7_2 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_7_3
+ dout_8 n_7_3 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdinv8
+ dout_8 out vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_8_0
+ out n_8_0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_8_1
+ out n_8_1 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_8_2
+ out n_8_2 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
Xdload_8_3
+ out n_8_3 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_18
.ENDS sram_1rw0r0w_32_1024_freepdk45_delay_chain

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pnand2_1
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Mpnand2_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_nmos1 Z B net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand2_nmos2 net1 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pnand2_1

* spice ptx M{0} {1} pmos_vtg m=10 w=0.865u l=0.05u pd=1.83u ps=1.83u as=0.11p ad=0.11p

* spice ptx M{0} {1} nmos_vtg m=10 w=0.28750000000000003u l=0.05u pd=0.68u ps=0.68u as=0.04p ad=0.04p

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pinv_15
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 32
Mpinv_pmos Z A vdd vdd pmos_vtg m=10 w=0.865u l=0.05u pd=1.83u ps=1.83u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=10 w=0.28750000000000003u l=0.05u pd=0.68u ps=0.68u as=0.04p ad=0.04p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pinv_15

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pdriver_4
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [32]
Xbuf_inv1
+ A Z vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_15
.ENDS sram_1rw0r0w_32_1024_freepdk45_pdriver_4

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pand3_1
+ A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 32
Xpand3_nand
+ A B C zb_int vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pnand3_0
Xpand3_inv
+ zb_int Z vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pdriver_4
.ENDS sram_1rw0r0w_32_1024_freepdk45_pand3_1

* spice ptx M{0} {1} pmos_vtg m=5 w=0.755u l=0.05u pd=1.61u ps=1.61u as=0.09p ad=0.09p

* spice ptx M{0} {1} nmos_vtg m=5 w=0.2525u l=0.05u pd=0.60u ps=0.60u as=0.03p ad=0.03p

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pinv_12
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 14
Mpinv_pmos Z A vdd vdd pmos_vtg m=5 w=0.755u l=0.05u pd=1.61u ps=1.61u as=0.09p ad=0.09p
Mpinv_nmos Z A gnd gnd nmos_vtg m=5 w=0.2525u l=0.05u pd=0.60u ps=0.60u as=0.03p ad=0.03p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pinv_12

* spice ptx M{0} {1} nmos_vtg m=13 w=0.29u l=0.05u pd=0.68u ps=0.68u as=0.04p ad=0.04p

* spice ptx M{0} {1} pmos_vtg m=13 w=0.8725u l=0.05u pd=1.85u ps=1.85u as=0.11p ad=0.11p

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pinv_13
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 42
Mpinv_pmos Z A vdd vdd pmos_vtg m=13 w=0.8725u l=0.05u pd=1.85u ps=1.85u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=13 w=0.29u l=0.05u pd=0.68u ps=0.68u as=0.04p ad=0.04p
.ENDS sram_1rw0r0w_32_1024_freepdk45_pinv_13

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_pdriver_2
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [14, 42]
Xbuf_inv1
+ A Zb1_int vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_12
Xbuf_inv2
+ Zb1_int Z vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_13
.ENDS sram_1rw0r0w_32_1024_freepdk45_pdriver_2

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_control_logic_rw
+ csb web clk rbl_bl s_en w_en p_en_bar wl_en clk_buf vdd gnd
* INPUT : csb 
* INPUT : web 
* INPUT : clk 
* INPUT : rbl_bl 
* OUTPUT: s_en 
* OUTPUT: w_en 
* OUTPUT: p_en_bar 
* OUTPUT: wl_en 
* OUTPUT: clk_buf 
* POWER : vdd 
* GROUND: gnd 
* num_rows: 128
* words_per_row: 8
* word_size 32
Xctrl_dffs
+ csb web cs_bar cs we_bar we clk_buf vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_dff_buf_array
Xclkbuf
+ clk clk_buf vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pdriver_1
Xinv_clk_bar
+ clk_buf clk_bar vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_2
Xand2_gated_clk_bar
+ clk_bar cs gated_clk_bar vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pand2
Xand2_gated_clk_buf
+ clk_buf cs gated_clk_buf vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pand2
Xbuf_wl_en
+ gated_clk_bar wl_en vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pdriver_2
Xrbl_bl_delay_inv
+ rbl_bl_delay rbl_bl_delay_bar vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pinv_2
Xw_en_and
+ we rbl_bl_delay_bar gated_clk_bar w_en vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pand3_0
Xbuf_s_en_and
+ rbl_bl_delay gated_clk_bar we_bar s_en vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pand3_1
Xdelay_chain
+ rbl_bl rbl_bl_delay vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_delay_chain
Xnand_p_en_bar
+ gated_clk_buf rbl_bl_delay p_en_bar_unbuf vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pnand2_1
Xbuf_p_en_bar
+ p_en_bar_unbuf p_en_bar vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_pdriver_5
.ENDS sram_1rw0r0w_32_1024_freepdk45_control_logic_rw

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_data_dff
+ din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10
+ din_11 din_12 din_13 din_14 din_15 din_16 din_17 din_18 din_19 din_20
+ din_21 din_22 din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30
+ din_31 dout_0 dout_1 dout_2 dout_3 dout_4 dout_5 dout_6 dout_7 dout_8
+ dout_9 dout_10 dout_11 dout_12 dout_13 dout_14 dout_15 dout_16 dout_17
+ dout_18 dout_19 dout_20 dout_21 dout_22 dout_23 dout_24 dout_25
+ dout_26 dout_27 dout_28 dout_29 dout_30 dout_31 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* INPUT : din_7 
* INPUT : din_8 
* INPUT : din_9 
* INPUT : din_10 
* INPUT : din_11 
* INPUT : din_12 
* INPUT : din_13 
* INPUT : din_14 
* INPUT : din_15 
* INPUT : din_16 
* INPUT : din_17 
* INPUT : din_18 
* INPUT : din_19 
* INPUT : din_20 
* INPUT : din_21 
* INPUT : din_22 
* INPUT : din_23 
* INPUT : din_24 
* INPUT : din_25 
* INPUT : din_26 
* INPUT : din_27 
* INPUT : din_28 
* INPUT : din_29 
* INPUT : din_30 
* INPUT : din_31 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* OUTPUT: dout_7 
* OUTPUT: dout_8 
* OUTPUT: dout_9 
* OUTPUT: dout_10 
* OUTPUT: dout_11 
* OUTPUT: dout_12 
* OUTPUT: dout_13 
* OUTPUT: dout_14 
* OUTPUT: dout_15 
* OUTPUT: dout_16 
* OUTPUT: dout_17 
* OUTPUT: dout_18 
* OUTPUT: dout_19 
* OUTPUT: dout_20 
* OUTPUT: dout_21 
* OUTPUT: dout_22 
* OUTPUT: dout_23 
* OUTPUT: dout_24 
* OUTPUT: dout_25 
* OUTPUT: dout_26 
* OUTPUT: dout_27 
* OUTPUT: dout_28 
* OUTPUT: dout_29 
* OUTPUT: dout_30 
* OUTPUT: dout_31 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 32
Xdff_r0_c0
+ din_0 dout_0 clk vdd gnd
+ dff
Xdff_r0_c1
+ din_1 dout_1 clk vdd gnd
+ dff
Xdff_r0_c2
+ din_2 dout_2 clk vdd gnd
+ dff
Xdff_r0_c3
+ din_3 dout_3 clk vdd gnd
+ dff
Xdff_r0_c4
+ din_4 dout_4 clk vdd gnd
+ dff
Xdff_r0_c5
+ din_5 dout_5 clk vdd gnd
+ dff
Xdff_r0_c6
+ din_6 dout_6 clk vdd gnd
+ dff
Xdff_r0_c7
+ din_7 dout_7 clk vdd gnd
+ dff
Xdff_r0_c8
+ din_8 dout_8 clk vdd gnd
+ dff
Xdff_r0_c9
+ din_9 dout_9 clk vdd gnd
+ dff
Xdff_r0_c10
+ din_10 dout_10 clk vdd gnd
+ dff
Xdff_r0_c11
+ din_11 dout_11 clk vdd gnd
+ dff
Xdff_r0_c12
+ din_12 dout_12 clk vdd gnd
+ dff
Xdff_r0_c13
+ din_13 dout_13 clk vdd gnd
+ dff
Xdff_r0_c14
+ din_14 dout_14 clk vdd gnd
+ dff
Xdff_r0_c15
+ din_15 dout_15 clk vdd gnd
+ dff
Xdff_r0_c16
+ din_16 dout_16 clk vdd gnd
+ dff
Xdff_r0_c17
+ din_17 dout_17 clk vdd gnd
+ dff
Xdff_r0_c18
+ din_18 dout_18 clk vdd gnd
+ dff
Xdff_r0_c19
+ din_19 dout_19 clk vdd gnd
+ dff
Xdff_r0_c20
+ din_20 dout_20 clk vdd gnd
+ dff
Xdff_r0_c21
+ din_21 dout_21 clk vdd gnd
+ dff
Xdff_r0_c22
+ din_22 dout_22 clk vdd gnd
+ dff
Xdff_r0_c23
+ din_23 dout_23 clk vdd gnd
+ dff
Xdff_r0_c24
+ din_24 dout_24 clk vdd gnd
+ dff
Xdff_r0_c25
+ din_25 dout_25 clk vdd gnd
+ dff
Xdff_r0_c26
+ din_26 dout_26 clk vdd gnd
+ dff
Xdff_r0_c27
+ din_27 dout_27 clk vdd gnd
+ dff
Xdff_r0_c28
+ din_28 dout_28 clk vdd gnd
+ dff
Xdff_r0_c29
+ din_29 dout_29 clk vdd gnd
+ dff
Xdff_r0_c30
+ din_30 dout_30 clk vdd gnd
+ dff
Xdff_r0_c31
+ din_31 dout_31 clk vdd gnd
+ dff
.ENDS sram_1rw0r0w_32_1024_freepdk45_data_dff

.SUBCKT sram_1rw0r0w_32_1024_freepdk45_row_addr_dff
+ din_0 din_1 din_2 din_3 din_4 din_5 din_6 dout_0 dout_1 dout_2 dout_3
+ dout_4 dout_5 dout_6 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 7 cols: 1
Xdff_r0_c0
+ din_0 dout_0 clk vdd gnd
+ dff
Xdff_r1_c0
+ din_1 dout_1 clk vdd gnd
+ dff
Xdff_r2_c0
+ din_2 dout_2 clk vdd gnd
+ dff
Xdff_r3_c0
+ din_3 dout_3 clk vdd gnd
+ dff
Xdff_r4_c0
+ din_4 dout_4 clk vdd gnd
+ dff
Xdff_r5_c0
+ din_5 dout_5 clk vdd gnd
+ dff
Xdff_r6_c0
+ din_6 dout_6 clk vdd gnd
+ dff
.ENDS sram_1rw0r0w_32_1024_freepdk45_row_addr_dff

.SUBCKT sram_1rw0r0w_32_1024_freepdk45
+ din0[0] din0[1] din0[2] din0[3] din0[4] din0[5] din0[6] din0[7]
+ din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15]
+ din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22]
+ din0[23] din0[24] din0[25] din0[26] din0[27] din0[28] din0[29]
+ din0[30] din0[31] addr0[0] addr0[1] addr0[2] addr0[3] addr0[4]
+ addr0[5] addr0[6] addr0[7] addr0[8] addr0[9] csb0 web0 clk0 dout0[0]
+ dout0[1] dout0[2] dout0[3] dout0[4] dout0[5] dout0[6] dout0[7]
+ dout0[8] dout0[9] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14]
+ dout0[15] dout0[16] dout0[17] dout0[18] dout0[19] dout0[20] dout0[21]
+ dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27] dout0[28]
+ dout0[29] dout0[30] dout0[31] vdd gnd
* INPUT : din0[0] 
* INPUT : din0[1] 
* INPUT : din0[2] 
* INPUT : din0[3] 
* INPUT : din0[4] 
* INPUT : din0[5] 
* INPUT : din0[6] 
* INPUT : din0[7] 
* INPUT : din0[8] 
* INPUT : din0[9] 
* INPUT : din0[10] 
* INPUT : din0[11] 
* INPUT : din0[12] 
* INPUT : din0[13] 
* INPUT : din0[14] 
* INPUT : din0[15] 
* INPUT : din0[16] 
* INPUT : din0[17] 
* INPUT : din0[18] 
* INPUT : din0[19] 
* INPUT : din0[20] 
* INPUT : din0[21] 
* INPUT : din0[22] 
* INPUT : din0[23] 
* INPUT : din0[24] 
* INPUT : din0[25] 
* INPUT : din0[26] 
* INPUT : din0[27] 
* INPUT : din0[28] 
* INPUT : din0[29] 
* INPUT : din0[30] 
* INPUT : din0[31] 
* INPUT : addr0[0] 
* INPUT : addr0[1] 
* INPUT : addr0[2] 
* INPUT : addr0[3] 
* INPUT : addr0[4] 
* INPUT : addr0[5] 
* INPUT : addr0[6] 
* INPUT : addr0[7] 
* INPUT : addr0[8] 
* INPUT : addr0[9] 
* INPUT : csb0 
* INPUT : web0 
* INPUT : clk0 
* OUTPUT: dout0[0] 
* OUTPUT: dout0[1] 
* OUTPUT: dout0[2] 
* OUTPUT: dout0[3] 
* OUTPUT: dout0[4] 
* OUTPUT: dout0[5] 
* OUTPUT: dout0[6] 
* OUTPUT: dout0[7] 
* OUTPUT: dout0[8] 
* OUTPUT: dout0[9] 
* OUTPUT: dout0[10] 
* OUTPUT: dout0[11] 
* OUTPUT: dout0[12] 
* OUTPUT: dout0[13] 
* OUTPUT: dout0[14] 
* OUTPUT: dout0[15] 
* OUTPUT: dout0[16] 
* OUTPUT: dout0[17] 
* OUTPUT: dout0[18] 
* OUTPUT: dout0[19] 
* OUTPUT: dout0[20] 
* OUTPUT: dout0[21] 
* OUTPUT: dout0[22] 
* OUTPUT: dout0[23] 
* OUTPUT: dout0[24] 
* OUTPUT: dout0[25] 
* OUTPUT: dout0[26] 
* OUTPUT: dout0[27] 
* OUTPUT: dout0[28] 
* OUTPUT: dout0[29] 
* OUTPUT: dout0[30] 
* OUTPUT: dout0[31] 
* POWER : vdd 
* GROUND: gnd 
Xbank0
+ dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5] dout0[6]
+ dout0[7] dout0[8] dout0[9] dout0[10] dout0[11] dout0[12] dout0[13]
+ dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19] dout0[20]
+ dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27]
+ dout0[28] dout0[29] dout0[30] dout0[31] rbl_bl0 bank_din0_0
+ bank_din0_1 bank_din0_2 bank_din0_3 bank_din0_4 bank_din0_5
+ bank_din0_6 bank_din0_7 bank_din0_8 bank_din0_9 bank_din0_10
+ bank_din0_11 bank_din0_12 bank_din0_13 bank_din0_14 bank_din0_15
+ bank_din0_16 bank_din0_17 bank_din0_18 bank_din0_19 bank_din0_20
+ bank_din0_21 bank_din0_22 bank_din0_23 bank_din0_24 bank_din0_25
+ bank_din0_26 bank_din0_27 bank_din0_28 bank_din0_29 bank_din0_30
+ bank_din0_31 a0_0 a0_1 a0_2 a0_3 a0_4 a0_5 a0_6 a0_7 a0_8 a0_9 s_en0
+ p_en_bar0 w_en0 wl_en0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_bank
Xcontrol0
+ csb0 web0 clk0 rbl_bl0 s_en0 w_en0 p_en_bar0 wl_en0 clk_buf0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_control_logic_rw
Xrow_address0
+ addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] addr0[8] addr0[9] a0_3
+ a0_4 a0_5 a0_6 a0_7 a0_8 a0_9 clk_buf0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_row_addr_dff
Xcol_address0
+ addr0[0] addr0[1] addr0[2] a0_0 a0_1 a0_2 clk_buf0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_col_addr_dff
Xdata_dff0
+ din0[0] din0[1] din0[2] din0[3] din0[4] din0[5] din0[6] din0[7]
+ din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15]
+ din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22]
+ din0[23] din0[24] din0[25] din0[26] din0[27] din0[28] din0[29]
+ din0[30] din0[31] bank_din0_0 bank_din0_1 bank_din0_2 bank_din0_3
+ bank_din0_4 bank_din0_5 bank_din0_6 bank_din0_7 bank_din0_8
+ bank_din0_9 bank_din0_10 bank_din0_11 bank_din0_12 bank_din0_13
+ bank_din0_14 bank_din0_15 bank_din0_16 bank_din0_17 bank_din0_18
+ bank_din0_19 bank_din0_20 bank_din0_21 bank_din0_22 bank_din0_23
+ bank_din0_24 bank_din0_25 bank_din0_26 bank_din0_27 bank_din0_28
+ bank_din0_29 bank_din0_30 bank_din0_31 clk_buf0 vdd gnd
+ sram_1rw0r0w_32_1024_freepdk45_data_dff
.ENDS sram_1rw0r0w_32_1024_freepdk45
